//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab04 Exercise		: Siamese Neural Network
//   Author     		: Jia-Yu Lee (maggie8905121@gmail.com)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2023-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME      70.0
`define SEED_NUMBER     28825
//`define SEED_NUMBER     28825252
`define PATTERN_NUMBER 5000

module PATTERN(
    //Output Port
    clk,
    rst_n,
    cg_en,
    in_valid,
    Img,
    Kernel,
	Weight,
    Opt,
    //Input Port
    out_valid,
    out
    );


`protected
+-94HJRc2S)A;X+8^R;fI7bHEET[Pd[=/PS/AbT)3JS[a_4SbY,>1)9IVAc[[>2U
[D,T+IFN>^>^:T@D\Sd.[]W/A)FC>#,)8c4@P@A<8<V=DB;(.8HA2XZ],ZB/NX-R
)a6G;DcN_QT<9M2S^_+9&g?)EA/@?gD74f@67c(RS6S7d&@R,]:Z?@YCe0K6eP]d
53MBJ<FNPA#R[WaPI0OfGg=RWQ0SRMCR=9(-e1;P=96c[P-YGZUfaL&^a_\4P]JN
c7FKd:^>V-\gTIK/^?WEMB+RdA07d9&()9BL_]ePEKSE^Lge=-VeaE&^K$
`endprotected
output          clk, rst_n, in_valid;
output  reg         cg_en;
output  [31:0]  Img;
output  [31:0]  Kernel;
output  [31:0]  Weight;
output  [ 1:0]  Opt;
input           out_valid;
input   [31:0]  out;


`protected
X3\\Y)I_g==^N,-JD,MDg+e0Q.TReL[c9.4^GaJg\M<40TKAbZ.Y&)&=GI-acd1_
e>MN0X6S)(P4@Nb=K:ML]DA0e/)aFBgRBFYYI<?(<3^G)19_,)&_S]V<9UVQ9::Y
E3b-eHBVc]4\#9c]G)4=^WK1TKI2JLdH+]F3[SK8cY@aVEENFF5Bc&d99?SLG1>c
NUV07:+P-;V\R.Y)_KE3O8[S(d)352,HNSCP23/A<aTTOASgdcHcW[5_e\YWR8eD
8Va#(G8]a(Q@T<G9,+.3\[-E0NdD1f_ORd74MMO_#Q1&-(3]-e/4DOO];UJTP+f[
-c@^1gZYW/He^J>J3QcLO1/@]eGWSU\JUUATAI6U@JCF&HDE_EQ96d9(/HDHFf5O
&FOI44O853O7)H]E2T-NCN<OG,V7446[B-O8H^V31@>RZ=#4/Z:T?__TC#CNB^]E
T01WLO?9#@,g.N\R/A+2Q&R5X9DTTg@SH7@&&>U48_W8KVPPg2E4+0K=UY05JD&d
aQd=MM)<)J89Tgb@A9^^6X[F;f/a74=)PF2IDBdI8X^4-f->c?+-^8A^T96d?O&H
?E&12(5O-<K]9R4a1F(Rg:_fIRUZX\V]?_\I\K04RY,PG#3VYM]DW9&f-F&b6Ea/
<1X78-]Y]RbRB?I+>Xg>fgM>F=YG]:EJ^IHM_2U#?YKV(01&;&;DW&<26N^g9Zff
:6f1CO;K3(),V+QJJLW@GDG4BgA\MO:-Z3SGaR92H-OcfRKK^M?S^F(B+IP>1_H4
0(aDLX(0<U>WRT.0>cI8[HBMYg,X26M@Z47#6<I/)WQDe>_B63<cZc+P/_DC<;df
W/=?VASZR]5N@eZ^ZJB\7a@I8@B=ND3&7&K:8G)?4:5b&dMCH]Q=]JLYbF,V/.:>
(DS83Q94ebdU?fM3?OO.1dB04G7EFSEX2@[@+Og:Le]]8N3L?JBdUXD<)FMZ]7If
gC66G-2a@DZW/,;03>^VGHTFQ)+0Q@:=b[48[<0_,.]VaQ0/2?2PJ(VI->.9fegR
83Mb:@OSBGSB54@]<.[8G__3a/<b3TJKMYfDcNQ&J)VM16=V&N>OJO7U>Qd7\C?X
Z^3>N>75cOTUa:db[+&T&(1SI0A2d>eL]^2QH33T(>^b6OEJa)6+eaFL;ePVCdB7
.OI9)\N^Re<d[0=>^TKZI.N9WG:XPO1M]C2eMfW:)C#(G?,70M,G@423+Q+cH3Pg
X),0<[38&G;^S1RZN2AED>7W7.<7DG3E@?:H8F(e-I=53.Ja)G,BA^DLGSbIEVf/
H-RBN<R\-MF9[5;+A7b=deLXOg=^a:4X&7?L-[bEN&G7cYTG@dSe_V:S>bdgKEM<
.DALA&V[MO>W6R-;NW/RY,b\]^-SNA5LL_bO-JLLc).6aM@.eL18XZMDf/Q.\dI&
[4JND(PR7RNb;+(gNASC:e;Jb[^4fY&&ENa)cOc,5?c#/@\DL4:4W[gGX#,M1JE_
bfD+EE&T@;-gRE315OL9RbBV?9W[,FE[N0-9+g[/+X,07OPR2+_ZaE[g9U4ScBR.
]D[L[TOBfc?5WGeg6LXP5aRc/^NER^c8RKD?77/[-UTAZ)6_^D+]7@#(]O3&&[R>
Q[N2+-&X83F^Aa4MVZe;a^U9PTAf;EK]Xa3(ab8V#X906U7[04;_\W;ZeETS3O+6
d?Ug,EN(eg.J-5_fLKZ]&WZdEg)[4\2]2(;a#-4Z.ZVRVHe0]9C.](7Q8N2V1;Ga
^90Q\VGYgYLQ))HWS\M:I#g>7=HPHGbBg-CR.dT9g+_e[gbQ^8Z&WKNOOeP(K-C2
IB;T8#eWT@-fGB/?M?X48DdKNMWZA8M^Za6bT)N21\AR<]C[17KHA6Q0gRYF^#F(
Ya72;#D+\&JMPUC)CJ3bEBe07e0Tf[,/+IRAgUW3G1V,#&&f\KO[bYCbN1QWY.C[
cCW33OKTeAg(0YTHQbU&9]<87?TZ;-fX_cS/\;LQ1LXgO&:G=Ib/P?QE80RefYN0
gPKKEKFQb5ZD2EURZAH--Ka:A/#3:OZ?]DHQ[YOX(-A?4IR[dc3QTL=SE2N,+aX]
cH4U5^8Rg]b[]]=bPHb]J;1)ASF-PN6P6BWcT=5fR5TFIQP/HS1TX81:(&D^@K3P
,<GS[D)LOBQF5R<gdSgf@aC;[7a7N?VL#N_NZPHP_17-eQE;1CMf]K89PX+gWZ-6
7?(D4;ggHHJ39D:f.:K=M][;d45>8HPOQX6,YXB:/JAW3=YOg-.\6#b-S]f<QgZ9
^Wc)Sd^?/,MeB:I7]ILD1c@H;@BU>>+,<TJ3@=FAKRYI=9\F4A>X@@>Vb-SJ7X(H
Q?CeS;Kd&LJX?Aa=eBEGV);MPXX=091XEa<#RK[M-@,[6_b\XLM+U9P.aaK+a.C;
7/^VT(fG?10[.(@cZeX1=+C[3I=15(^NBb@3:VYOD=8:N3F>1?@<8Fc&^3LeZ)-Q
D-_gIJDUN9C80[KW)@3Ae6)0/\[9f^fJ[W8<MEg3#K]@a1a).N-I[5+#1XAc8RJP
C3AYg40;Uc5WE<SGfgI-1KMC#JB>\1a_H#YDM)UZf(1bJSU3f_GFV]&f1eM?Q<XE
d(8F<e;Q^aEK4>;6D73=H8PLf[RDWa8gCNA_WY+2A@V-17gO)YO\A?1;d#+L#SI#
)a7E^R>Z#16BeO/,O@)]R#>a[5^7P/\TK8a7,RF),cF5^1MJ?4HI328We8/We\[9
=-&?d_2a^a2#cLMf=M+.S^EVbTL/S:8#+O:ZSP>R7]G?C>H&a)3/cR8B>F:4B/-c
=9F&<:3Z/=.A7C^_X5^C,G,.DcL)+Xgce6.6VM,(ALPQg3&=S5/&0O-N9[T_Y-^8
-U)[]E9YS2-_+5(QUUO0Xab</e<G=3E.Q=IZ110AC.KYJ?H\9.Ze5P4@Z9)ITMfZ
UT10BU++NCJ]ZL]K6E76_<>-A>IL;=TWRR099LeO;?&[#B3e4MCS-&dF-)QCGK_,
dW.KMHW?7BYc6?]/>Kafe+=>Y#3U2.4)\<<.eZ+6dfVIRPMVbLCe^42J?;D>&Ua2
3\)(g6O-A1LYJSCP41?7?_(04U_SfK;_3cdHU^:37-75UAFBAR+6N#ZBeXZ=I#1_
B@:37_^?6:d3<^L6_B)(eB]f29(>\M#4fX;6BQf01\Y\KIPZD>K+HD0\c.a6f2K=
X-+9J89TH?ML>_QN.5\-Gc22_AACX.Rd-L3P@LeFf5YG&UOaDZeU#=BBNV]GAb(^
9Q^.0C6H:/&F&XXM<1/)3;R;L0I:C]fOTU+aOP?+dWJe7gZV9670I25aOJ68CVe[
5&2^gMHJ?gb=+M2\C(9VY(JfN8aY_15?L)I^>/<HYR>#3?VF6<?bE.58EBT5U7<H
e,OafX@69.e6?<_+DSD1<^^YV#eb_gCVdc?DcDF3I&,BFN1g3WN^>?ST/)DaX+#&
Oa6-15XEV?QYFOIF-Z>e27-D7S0KKQ#JgJC=ZC+XQ19d\&;e)U;9;AZPJC595:^E
ZB<cL11b<(GB\.WG)M=Y[G.WCcHa(8K3EA)FLEK,]45:2eCdDRO7^N7@eV23ga_E
GdJ0V@Ccb)3?8E=)_=NbH-<GNDDYQ>g>EbJbdN+BfWFHH(^3\3Pf2+&S,b]5V66J
Cf+#]E^]Lc<)2RQ&X]J^I2DA?J50#5+2b10O-JW=+a0GS_K31I/U<ONS.R_N61[J
Kd6G9^5YN)E&;A(XNf37fReYT2)b_8P\6D&+T>M=,G4Nac<GVdP;D]@gL>@FDd4D
]UE#KUF@IObL9;dY#(M0D]Q=cWPM8fPG]@0g]#_905^#T\=3J^][W<#07:DgeaD^
6Pb:dQN(EMNc[E&98g<XU:B6@;^_-(aW)6V&0GgZHPg<3#B0X)\/(JRe3.Ub-^M<
)2G\J@:b-?^6^#=#?dG54[PV+_HX\H6,b(M2\?DS5[CT]#KO9IbY\UA/TMV<[H.g
U(<41PG-YK11Kc[DZ7#T)L9]P+@P(b74V.ZT\:W6?-b:7WN_G0)>.eAY[ABER+S#
dOT6I2.UM+^[I^,LP=,I0^X@L^a4609^=S&Y1_a#dE\BLVb@I9^7?MdGB0&GKD@@
b:5]S0.V<TY^0?W6Ya(Z:F-e;\e,3bDK0OK]64XPa[f)K@#^KG:EN-]EK//[-W+c
QM[EEE&4CIOWQ<0L)W=YIc+10UU(#DYMTY;N(GGb]CZF//Ta^9)HT9_GR\=)]C:/
EV=4gDW=<I#aAR,IKU@;5Z.YR]6,.O1#(&4Q@&V1gEY6/b38>^_/Cd5]IBf\@5b/
/7Kb#=T.]LT60S1UBKF?01?-2XB1[IR.a;0_&gbGdY0de.TF84V0dXc#NDJ..JKC
P-8>X;@_L@DDa;WKG-^,Z0/CMV=d)6J>d[J1d)LQ[=#ddc([U9=G91PZXSVQ>LbS
7.1CA?09[6WfQ#Dd7b]6@)\+V.LB&\@DUL+P-4OWR^=Z_++FXQ)8LHZZB=FT,&_<
EgVWOOb3]b23[6BTc=8/1]NHR+c<ec1M#Va8GB\\I)A.@HO1cae<;,9)deBaQT<T
Xa7fNH/8F@VJ0_:IY.;gY3L1QfEB]E2)Lf,F\ObE(bDPHB=,/NWc7f#W4CT2,Z;G
.4C-]6bC@N)JYV,.A?5gLeC+[8?RBKWYV]XaBeRgOF9<X56YgVIO+^+f1H[VD;-)
U;f=P?[XaGL@5LFQF[Ec?00>Cb==PNH)BaQON,\GAa]&0T&Y>OZC(.V=d@,.A=S^
UL2)f?#(A##N^^3,d)^.KJ,=cGDMe:Y:S]JR<JPM<O6^^OIK@IG4DM//WLJ9]U)_
[(9&T5?^9@Cd+L7&P-NR<:4O]JONH]#K50)b]YG>JBUT5f6(.Aa5&3:^.UKY([/B
:RU/+V4EZ?a@8CW>2^V-A&VE;B;G<GeGbY=)c=RL?GfAM_R,HS(T5RUT7H9LADKC
2>QO(4.N:#[77P79TYgDGV_I@\1.LC89]@N,5\\gBCg8>M+aSeZcFO;KE?Z_<J3F
?FHZ9J-SV?W5)YZ@:2gW9fR0\J_=dV50&@-3Qd+7T[_MWcRMEZ/)9SbL<QAcC\0K
+G0I79&8W?&OH9Za:9T#\9e2_S,&J6<^#&K(0(<>WHEK\S61#6SJ#gRF=b_^gW+_
Mc#f?L/832;FDa>G^]J#,_7N,TYKK1R5^/F-b#&S8(C8G>,=Bf;TW=L8<.Y;(PPf
ZF6_4?bKO)e)b/BZ+aC9C4@6;+T0Q&Eb7:V+=G/Cg7&#a]2F8G;C2bC?Q51e6^@9
==EU@JA[MMHMB9AXfGCPDF2<.T[5e:Ue&=1VKQ_B@@D7-eG;>;/Raf6O+TUP:e9K
G]<C:O@/L59+VJK@PJeVdV81VHSc/d#^&[X1d?a9f&)2JE?O[KDWLL3cfD[2OI8O
#eC-b;OB_5g<7[N:GbA5+3b\7CCa_,^+bY49KW0C,=UV<gM37DM4?WDTL+PUR^]M
0ZA_#D@.W^IeG&M&X\AWZ\:T)C_4Kf\fLX4dGc17Z&UNZJaCKMZc7)>U5:PKW]QO
SSOI;b)?@88\E=F9Q86R6L-0ZGK-<(=ddbV(J/9.V=J4-3^[XQXgcB4ZRD\9W;Kg
#5;QE:D8_cUf8Z>GcJC;X/e;9Ke(b7E[-8^&\:][;3R4D;=YV/ZCf48<YQXbLLU.
2a1#T72^KB9_OZbaMYRd0AdcH>>_XAeN7a[VE,<MY5PD[?O^b.EUQ.<2Q;EO9VKM
ebA:,DRbLV3cK(VB04Y-WG1<f\:@609>=.4Nb6e=0b[g.OMEO4../3MR)/d)7ePP
GG=<6G6afT3P4Fd1ZEbJHTAb#0<GVBPJV+d.Mc/YTgM0FST#B3?FSH?;AV+NQ)>R
:6DK#IT-^JcJ_OU>8DH^5-b^R<IVAcfG;VaM7M66DH]-X)D#H4.>M_[:(>8E3H77
0&812=:<+]0HTTIUU[JDW&<H;KNJ(R6_8&UAe[Jfde/PWO6R]=2a[NL_@HP:+-?#
3Hb[KL#+<TbP#NPe2FH(gVB@;c(DVZF&9&2Z7C8/(M&<(cZ]UGWC=PB\;&O0,a/F
6DD8;cTGeR8;41fU^D6b0?P/<GBf#T@g(M&,,H42bG5bH2JCAM/\C8M_[C&77K^E
c3\&+W3>A4N-K4g&S7d^a:Pe^/V2XAa7KV1X@GCRaO>3:H?,9KNCI9fFL&c,2:1>
0&IA2e\AZKgdaYTUI+bIAHOY4\5:M__JYUd)D/=a=)QCI6+@0BdLY85EaW3AXfKe
]BC<,?L6\O&^W]?#T](K68g6OWR_WCV_e?aL?_LPFGg>(b_Z@J1@]3O\D:J]3PL.
H,\/afc)N,PgH=I@\9UW)8H/]f5XQS/-FCZ+1HJ<I?d5fD8fU(gV_8d?1U,&VKg1
-^Afg>,cA2A/Q<ZJX0>)73BWF,.W\5T]GQ(T^=eBb-QL;T?&-QJVAII<4d;Q\L<g
63U<4L5D[23FX:d.d8ccA4B[=feR>SQg/+AE=e-a1^@:(E=6I9>Y+aCEA,Zf#8]4
<cB\H2G/;&ICZN&MP_1]I6_C9f4FXPaZK-AMBFUWJZX]?24;H-I[JcGQ@:N[+-MG
.O#/2LB57VECK_DC^A+@B3E8@](24UM\/--98B,b(<PXYE-.0>>\UJ9R[ILY9\,<
:ec[[3?C]Z6S-3>TFaTD.9TAM[ZZ44F+YIG(NH?ZgY,efY]Yc9G#3&)4a2[7/-f[
Z&X;,<P;PYXcf5:6)cXd/1=a&6LXQ4^T>g;).H1d0/#:8:KfPa\;)0P.D.DUHFD/
=R8Nf>6FZGSf>ZG<YSM@25JMHBaMH)G#&50bU=Q@5b[1D4U5_g_F->/B.S#P[@^O
ZeB&#=GDJ45OEce]-g0]9\M?.?CaCK2&YJ<L,ZAg@KbVUZJC][IZ3N5gW)Q,_X7)
RBG&b(=YU&U)T<0P_e#0)B:1X860=,=AB8PTWe0J/#9fW1,E]9)+V&G.+#SC45aJ
SYWCF:U1Y8B4MGa=/ZM--ZdFY\ZJc1:c\Yg6ZTSW;BD86PdE8D@d6R7U\K#5BD)P
bG)T&Z+HeAU:Pe)9H+@4OOA0d4SQW[b.=/5_T:(F^_3<JIa7LFDQ5,fF5A(&c(JF
X@\C^,X8:,>Y\d0Y24&Q#J6:I1.EeTM30ADNN0WJ9B]/,3?.:G&[MOA^6\-)/CQc
+2^PKbC)TPM0G9D@YdF>ae.83D.<LW.8g/X3/ZGUZZ28ECOH@EK9XB_4]@E-?f.R
765(:(P03_U-K==2g/TCU=B\c8W7;+KR;BDG9g7?(#E,0d0L66:HCZD(QP#)?5@_
ZeTQQfNFRMXP]/6K-?c(E;#bd7N43Y+T4BFL,4G[?&]?LPbNL/H8YDS&CF.Hc)c.
J-[3Tg1QJ_[9G=/5+[PORDFMT-G[<[/f4I9<+&_;2_:Qf\a?@69fJ)GPA]=aJA>c
^,XE2Y0\-J(Td6)981>_:Qd7P_\H=[R<4Ff:cQ7M]].KEe78621TaMcK-DBLA:f5
Hd)EgKN^U-f,Ka\[DdB=8.\#/..#dg2&8JNJ&R,YK7:>)g8S_A=SA[L42+42G0H)
,8QGBR+.K<1a@JA.c;NE4O8b[R;Z=2\fEG4.<D.T>6>b&69JYWT1+EFcD/aGU=C&
=/2MN?.eBQMC3#a64HKA^NEA]55G7:.]\:+3Q@(0H7X=&P:AWD)]9MD6UC]cIS_e
e(E_ac]E,5/2c&1EXbWG)RO:cF0J+D-?)4_@(8-a[P1[^[Y#-g3R2Qb8Ie0O7][=
RE#H2.&f.UC\6f7AD+T74Y.gA)Q@^@1Y>YD;-:3D^]0gdS&6,:1c3CX-1b(e0AF1
&U_;OD6FK[1CCUFIEWNF2IG-/N,9,/c7CY.<<N1@/#[7G+#S5VKcRM#:X__ZHO-P
b9=D59I=3G,0Ag92-(DdGJKCS&(L2e47K->bJGfe9X2SW-:#A36SH4S(4eXEDcPN
f1ge#b[>A+\GZQYQ4&b@[.FSNYG<22QY=ec:W^/YM<J[HQ/RfZQZQZ?C99\RNW]V
:UK<bC0-BE_FOS\L<g5A8W&]Q.U3XBL88P2Y+(9#QV71O6,N?RC+/#-=O</^\0gY
?IaP.0H(&/H^]@MONFEQ1T0A(PBN+(#R(8L@QU)Mg;[_/D8G9DLe]9UP10A30]0)
8TAQD@29PEYM;&dQ]SKO[E?D;7^8R?V1YR<F\=0@-OeW:NCg_@8B5)/g1;.<9FfR
=L6FW0CW4\9g0T63cTN=IB<,&bd.GPf=7YIC=5gN?FDdY&[()3R\fVU(X=HN1,Rg
H\3S+8)&.L7H7c>GG1HW4(HA\@W[:.=B4DY<-O&H9M4GbbN=2[_:UV>,a&Q#:;A(
XfWRM2:aQ6-[94:D?(R^0#KKX)_B2;MB/7OVJ,G2=Bafc<;9dgNOHQARG#aVH=:.
Lb0dMVIPEC,.:YC0ACB2]=&IL.=_Ee7g<D3>I10MK#HU0_MZ3W6DZIf@]BE#<#3W
:0S00-Q&/O-(b#^[3CUT8F;RJEA+b8c#H06&.XfUIgDKG#SI,P\_M=X)]Zf)5M9W
/3LR8A:U,_6)?O6bL-HS60aBAZO#&4(S&&W7@&ES.S5?6)]^?CYXXKCMIU65^+EH
0-[\(d?=MAPgQUFS-EgaRL3\X<W6]=Fag?4L;AMP-KF4A(C#/Eb56B/R+4U_/bG7
cM[[TfaSQW>cZ<_=>&8M&J_\.CDD[V]=C5UC(,Qc:SM-TgOUK<1Y?aJ@7Q88>M8E
0OY,#f]3Z1)Q#9U^:OfE>7N/W,2:WS=XeD6UER:E[@Zg6&S^R?K\e@UbSZVgUR6Q
b1J(4GZXEC^5)I-48eOXX4CBL,VY\MD15W?W<a7,#AUNdK?)8P=^/G@bPVM)&WdW
cGM>\0f\dURDKO[SXf1eJ)/@\c;OY8dE<?MD+6?Z-5[02^eJNO6)-U/;]a3O9^bd
FJ83^OBXY+8XgJNGO[R@;cI4LFE/(_&@+&OIYc&-Ad:BCg^?e<H5_UCGd(0INbV\
(&+1-95:45C_1W95M[2]/[<QZ77O,<VA]XU1/9=f,UO-.Q1U,2A/J,V,adb1-GNM
:_TF7[#^>Mb/ZMM&<5&Ja^L7X-S0N_6UHQ9EPRVEQ9Pb2I,K]ONQ5M8>=K&=a&)/
[SV;O<NEcH\gMMZOIMUGG^Z/2Y?2>29DL5f7,S@>P,;<b]Oa+9QK^15@#K<5G3XH
KGgY]:8-;JY9T8?eU0O=JJW0/#A54f?HZYdC,Ff.OJ3C<][@<Ag(bF8>_J>>2D8W
a8EfDaWKNc[ZaYH(OI;(V^F[64I+I=0LH@FG>e14BQO.f3K#NZ7JFT(-:.2g3dOZ
]LH3Ra47+)UNT_gdM/J2>5SP#KF5?33@\MgE4afL]RdbZIM\aO)+cL7(=ce+Re?^
]Y,>::U2+BfSe=#,HVB99-_eOTUe0A8F2g2Z/EaAGN25[8A=W:U4/&(?F3)EN(]-
b]<<0+MZ-LaE5.5SSJf0-A/a?G.6LG_FI?+dGUCgH6^B&4]-aA(IJ9G^);[Q)5/8
,a8^e6c/I^ND]<HPJ>EP(ICZM2cc;a[a)B<Ig:;.9-_J5+8Y].(74YZ1/1C_T2K>
X@E2^63S)/GDLe;#<b6dY5MATI3[Y;fY9O89N=,WXO+KM:SCJ(EMGS4E[HS^9TDH
P.0DC:9\cZ_RJ2&-[+d_O9NZB5Q^G4Q5=1eYe)NKQFe;MfeIT(.._XNUBNQL>60L
fLIF3BPeDQb;[(dU[SEKb&U.gM7L3+TP5;ERU1aMVa&B9<YW/C+W2:TdAGEG@F2V
O7FVcQE+(M/R7/NZ-DK4Oa<[W^.J[3_YKf5(C)0,XHW>QGa^73Xf0DYIaQ5D;c&G
GK>(fX#&7Sgg=I,ADI#_gb>NNFBH0\),gE)/UCB<Uf.;-+dg;9UFTW]:O4\/dR@6
d9#G.+DN:H+#8=@.>3/R+APb<M.SUBTY)d-NMD=^Pb.;S^)1_]>PH]T,^^9=[C/e
ZePaD4(QSfdgAA4URM==R.1L9]G(@3^=aWfE-03A4SMbDJ/fS[&LNHd6?>MS5gGC
WYA>S,0LM?B;(TO>.6K;SW7FcA.4>fUR\T)@IVe<H:W,<LB;;#;fBO\JFGW,55=3
/7^JfE(^4ZRY<7+J[_.<bK&6[7OEKH8V[/3Ud;MeKGRG]]PP1B[(K8A?B7Nf[>d6
/Q-dAD1@(0(@8]K^Q>N+f7AU#RYe)/cRQPCX9-Je&<^_<1&V7Z_aD.(R()TBU5H/
4\]W-FN&)/Q#U@0a#;9^dT_(c6@?aZ[[;PZ@.Of&.a-]<CO.]9RSAdJXU-]+;;#/
bIS#d,c7b>Q_)7:(:,6Q>ACgPb\6A6&^H9.C7M;(Q7USI>8[ET)]Q2EGKf&>&XbZ
[P,6N>>0Q(.UP9=9)XMRH1\PLB<.Z0J^@:Q9GD<W,:)d<Bb)[C(cfDBNL-P4K0Z2
W:c<+CDDJ)fTQSYS]@.88R\)(QCJ+<LEPcPc5B_6^G2-NPBAXXWK(M/[.QA>J&#]
L8.Iad1,V+/7_+TYX0NEUX[7E=0/[[Yc3A?4;e)dC_Q6O8WfGP5>M^:QE#_ROc9+
Oa&:7@cQ5GQa#4+^d&5.5eBYS\OB4LB[VF6g>77;4_ScINWIU,d[#H3K)L;8U+XA
T-1a92-bg>X;_E>&E8#YBCRb?/8eBg?Y,SJGC1C=1b=bDQc3deJf2Q7[112?1Y(1
WQD&;S^>MZScg\a5QU+\EOb?dE;DY6K4aY2@eC0-N,9:PMJUQ4_0HA^-g<40\?#Q
@,Hg.d+adE9;2F)PVK(Sg&+O_D1I=FVV=\O^^R39W?SOA@T,5b;.)TE2=MNLTZQ_
,45cM+57Z&IK6)36>Z+XRD@)g\DJ&B3)+a/&V88:ZZ>FF]+/:]V)aX:)GDG_0CS]
,/0c,XKNV(2f6e]bU5eYNg-K]/5L.>:5_AY2LWI9G;6NA\NR6Q.WHR76T.R+5D<O
R/:G2f//C_c7faHKb\f=ZIT+QgBad9e\gSEF1S++IM;b7I<RTK</fALYTg3/#aLH
CH85(U&G[M@N5T_Q.:a<]0&4>P,.VNH[8L6:4S=,8bQ1W84:_A#d+4@[6If5U\I&
g)F,68c,1B)cIE+a#R;^d/0WK3Yg3Z7Lf>1L,CbQ^\CWGI:J0O@3N2?UgUX#a#f0
fc>-P37/A.HC3@PLR7T.+9@B9\OB_<W;O##5U\:6J\9JQ9FEeHI3^&dSTJ+;Y&TD
U\U<[6aI^5))a8C9@CIb(N4SU,M&fZ[=^[4-?::7AcUCK==#W[APO>=U8YXJg)\0
,.:bE@D=0P8V[QdJ@3=QZ[I?:K9ABGEB[M<#.<8JMRFR6,AK[aI:(T].OGMBTNEb
>Z4I+O\K#/O\EaGPY1J1d1K)/<=I,V;W@;:W2UV+WP0>(Q1\a5-8@-VXfP=WHI7/
KEZ(JS>>SSID9cJKf_F8-?\R=377LL^>,C4PQKB17I?Y,fK_OQ_N\\P9.(NACKF;
a^RV9MT&O[>K37,Da5MFO5XY,745&R,EMPR3)[DY9OdbHCUWe-\V]XX+FR76(/L^
^2BH\V\0_b-UR^I2CA9KS3QE5TIWX>8a,Cb4?0c<d?MH-R;@S<M?PaR6UY44.C-B
N)1\RT6<b\aG6TG6^M2J41Pg-<OSXf=_>cGRge/Ye#GIA(#G&K9NWI;PMKCLX4=K
]HQ4U,f8DH.CUCd))/=6Q+bDLS&/^O+P-(&IQJD4[M4//cf#6I/F0NMd.3IA-_3A
T9fXd)@YSY^O>6MGD5[@e9_N=W-:Y7WH-R1g)^0eTB78U6Z(;eL<8Ja^Z,O\OK=V
CU\YRB/^7c,:)K\4+L<T:9b&LYGHYHW5FA]?ZA^0/e]Kc-?Z=PI-PMK2>]43XU^I
#VRP<<)34Q@^4D8-Fd6QJAJ70<3U=]g?L&ML?H?bA[A5bN:#8Ga_gJ;(;/0/[9AW
H47c?[6>E9-fPGM73ZIV/CNB4A9]_JJB)97Z^[a,aD?E=G>,(-3L,[)_47N&PZ(@
R,6Y:[P5_E0Gd#Z;PRbK,IE15.WR41MYLgA.g(L1W-Q:41>/=EJQNU@M4J4^<>F2
^ZJg@IVHJB9]WTP5Q=],L&642f\T;JQ]4GgU0b>RZRPKRTgO^YRcSLb3<NQ\T.JF
[^#3TG4a]L.ANRKHf7C&cG^.0KIS8&dLWd@73JSO0B)-8WUc:;+6-RgA=F[e[Q6-
-BNRCY=9)ce9[W+dYa?EOca6IO^Ea/ZM2-,-N1e:.UICBJ/fN4A7^3MTO5gNTZ\#
XK6b.(_[JU)2Ye/XbTY&RT?Y#&9VRG(TdXQFS-2O-b,I&];934>NYW9Q\59=7fX<
0FYM2S,SVV;[5P3;3V.90(?M/3;&cc2BMNM32.S#9L/ES4U0N[[Y8[Zd-]^D<CH1
d<Ad_3Sc8>@5^a#)?M5:^V]/\Ld77gOM=Z]X6@c-f\FBZ6.@9>8BSU2#1:1aUD0&
&-AT..YTDZ&4ZRd60(::Y;cFGMY+Pa(50C7.D@=V6&R5S)e:5AK.>Z4FbC12#1,3
c.>NedHT20[)Vg50EOT_3.<7@QEDeP&W)ZU[E#V-3:H1OeNa7L@[>>48e\?A-2V-
=g4\6?WV=VS^=-XR/9U&[XGKB?DY8S[S^-?@b_VND]c?,E@c(I83SaP[e3bE.BNH
:-YegAc^^S33QS<>V4a?X+6\82>+VfGf\IZ:/b5.1\/+E0Zb/P8>+cF[@S(<b+OO
[79UZ]MeB&eI\Cd0CL^2@9,K=<D07]+MIBTdJ=.)J7I=B&H^Qg&HN75A&G\;ZKa4
G4BK:&8#eP8AfYOgeXBK-/A(<XgSb#YL+KI]UPEe[=LMBE++UUG=XEY_2#N^H-J.
<WSS6;_P)4S7ZaI5B>M#BBg;Z;#YP6W]a1&T;@XC).V[=N2gE:]R[f@Q,V&T<FGW
W@ZH:?+-/0dNMc+78(O2>/9?/fV>7L,<4A,BS]BSWP_IJ)abP]:.8\F&TBI>DgEV
G+\-X+1;65XN:I/39H<_S=LS+0.PAR<8L;BM>7g31F_AeIJ0F;EO)Z#-(g/2A@GO
-fG?+SW-9:6OCD<4Y<NWI7^2g19DG=(UX4gXM:PU5S(_+F<,>OMQZ[5VX1,d(f+M
Ra[.Mbg3.Z6K3ZIF[&\X>=ZVMJ,;e.d_cc8Xc:g_9R:UD)UfD\KF[C2LR.@4J+#+
Y./GK[8+:1WH=,d<C5H+V&-Y,[5?,CI0(EPbcfbCN1LP2OSPM,)@4e:==U;=5?D<
8L]_E87;Y5E2/&.:gVcK>@[]:))8WPZ[ZPIb@UgbL.AJM-DMZ7gO+,6]bL#C46L7
<fYP#fBe[b9>(ZfWA<@C.a?3>TNTK/G#AE)W1K3:6Ke8GZI8:SS6Kd+LPPS>IP]b
F:4=.^a_<8M@NQ>]Z4W6W:3U_-559@(R+?&1TaWF.SI&:E3.ddbPH-?D9dcgE7aB
0Y.L18A^\&_=00KR\>bW.\YO^#M;+/XHY^.<?&b.?L#Q>ASdT#7^L7TZ((^S12Pd
#O30bB_/(e<<S:O/1U..R#J17:2UFPdXX&:_bba#<6.#07f5I;IaOG7;d+aEO&1=
4CFO6g_GB>d;cf2S5>H&NT3E<V3AAGb7EeJ5gbVL2,6CK/(#(QF+]61:^6=BI[Ag
&YXAVf)@OI4V,&cO3AD7?f8W[0FN+7g^_Xd,FObO=4FI\f:ADdCg#X@@PJ\ZFgCF
A[3Ja&4b]-8UY:HCS/,.V->H66C_:L&SQa1L:-=a#\6-b7(=#Q2?G<EFT@#>S\8Y
JA=NOR<P8<:[57X7&B;6?Ff[S.YbK_\)VET.H,QX3PTa[5)/QN>/W,XJF[c9feDf
e=ObW\I2IM:HU\LAe]SC28J\&GL(IJ9968C6VRBC,F36N)T\BfWBD>J9C@E=;MH8
A=KQ2g7Y<6M<#Z?9G]5QF(F;]CA.25MT?M+LIV=9?P.cKM_S.C/ZI.?W=C3edQC,
]QZV6Q(ZGb;f,PLI];4=D<W,bUYTMK9SP/YW_4SB<B5E2Gf4CSbfMLb.G@PTgK@b
,#.T2ZT+M04&I@4Wg,ZZ>A\GA1;]9/CU52#dK]4?<>@OR;(CT,a_@.N2YQ8;a<9]
D>:B/JWQ?U_K+#IVP/ENK+H]If+3Qdd[;6B2<MZWY7UdGf13F5\+_cOMM-?,J/(^
H1ANDFAT_+_C.+7)K22=C,XRbNIQ7ON>_D2G;CLH8EbA&&bINX,;=b4T2cZG\G3A
PH_<BR1>G;+1AE5T9P+(EBV6/_9F+f]6IPf1=(V,^2V>U>L/+2GgW^_YX-TcRNdW
P6C]_d5U6FW6gSXQU4.?VVB)MU&b3;_O.NBWY.P=?f9[IIP\X+HG7[/4W?cJ]];Z
RM_:7S=bJ;A<VKW/f-92X#Gg@eYf@(V^;)CaD/<99;>E\DSHT<R1)3S[T(&^-&)>
gU2bLIOeMbEHA4B9R@O8G+ZVfJD.&@JG3a8c26T_ZGFRBd(KMGUELP:^IA8PEBI]
4(N,;YWLW8BBe2DJ88Z4>.IQYAY]6MW(+EH-bfbS85GC>DGEg)IDa=W+/[e9V\1>
L>WQG1=68FW0=U5Yc[U+d2<U^^G=J>Wa=[KdWd\7bWHCL^S:#^KB21V/E?X.>>JI
X+H/W5U_.3,;WEI\EL[0^9PSD@WbZ8Z79LJCGT5A@D<(a8bBJ2B@T:RS\A-?_Q@?
,35,<Y2Q(O@=2C,74(JH88_0]5GB+TX90R(7e,:07WHP61eS]ENZF/4;51<@QN@+
9\Lb.?I&HW49<05&K(d41QdbD/5&IFPHP2>CaDI??(4@H:UO_VBDJ>f,\6GQ/0OO
AK,&+9T4,JWM>;K-+eYc+a7/\?^ELb9Z;D_[A9Ib)PA>UA[3ITVD\X^Z=;,SO(/X
VYVdJI&CI;&B^5;J>8KGC#XR.M-?YY7,:E+3c^Vad&7R3::]Jb0M<f]CUA;+#6C2
/E#:QA7[V-(f?G#ZH\aM<R+<NQb@FeQX=FI,<c&bKNV?-WPVM^TX2FJ,Sd[A^OJK
AC)(MffE.R#7A55(#HZaLM5M#F/;6G3)4(<,OGYb>JdY/S2HY_6aAV>Ua>e(1U<X
MKW2:Id_^TX;QXLE2>d.A+[e@,2\;f_R0YdW<S3?1H+KJO8gc?>,#<8JD@E]c\FX
-Ce],#IDfY@)76B:Ie)6>dc@NTQWSFR@SeT81_^5-]c.-2WXR_0(L^G=H6FTYYV)
+bIeSZX].c4T36e022,e2]Mc1IgM0)AOI.ZZP9A^073<O(B88(H>+L4KC[AKg;bX
3ZaMcbb3PART9RB[G,A8\b2[A@R\JMN+03T3:5T/AZ.?IQC4=;IC/4P)AW1X?X72
ZN]I1X\9):@c#2=c2g_#U6QAXSC=<X&0<?=D\:ZcXDL.8T\(aDYQG@A8eAQL?a4S
VD@ffXP5e/Bb;dcG<-?VC+HQVF[e#/BTHMM32[4M/G]H^a]2\U3(H:D:+E3d)UTY
?.eY_e,KANKdL5HR8C?6YJDO7e\[DA3:-b^aIZ>^.cd(J,a,;GOIU-+@FJRa@KKV
],XMA/1)EBZKLFDM-a>[G;>)#V12.;VY2MP1=V+Ja6/^L(d/2feDD].fYaE&(>)I
,b)Y^95L5_OMDDOaE&gg_UHV.c^P4e20M:3:+c;D<ZI#ZX&#<UI+UR[/B#[,aTPb
3(+]@&g&P]f7EN4^=\E.bW@e&LYQS1e4cUO<42XYA4MX5EV\F<P>6;QgSfMSJPg1
S9J8d.LJBTDM<0B.J6:#@DK-7\ZZXD@#JR4a;#NJ+_LN99]P1U@[PUQ7EDCK#:A1
B>8cM.EbL7Q^1dIG/dQ3ZP=bCU<\8\R.>I[O9BF?W_=(KHQD3PSDRL4-/+,R[,<K
ee=#\WZGGN>-JLFI=/JG,0/T9NFL/W;+;#;?a:N.W.AIeD>:U1\PS:ET;_0+e1Se
SNU&,RZ\8[,CCQBg@XO>(3_X^94OVV-8R632e.#X5e\H&N9F]C)aDQ-&P66:f71#
P-RPZ1K^E#,Qa0WGaI+VBHO5@FWd.:+S+g;O[H&2(XPS-D(1F^\BadbROFD6Q(LE
g:K45Y_Z+6Y>CET#,A-;UPHEOcSJQ]\]?+ZQZ@U=<#,ec>O,-\Q^R/cR)<@^+FUa
A.JfY#B2R\dX[7/5OJ_#6-4F)-LY0+1B67dKU2R]<,-g<dDD<DH_)=63NU\_&8/Q
(WN4bJBSSW4#TdW\gT-Q@_SUP1<DJ)J<>ZV@_3:7Df4-c7DE.<J:Y0YY(/I?3UQd
F0?SAgOfPf0eR4B+@IO4B_g,K.M29F7f-e<2&CC)WN2WKVMJ#)V5,D=A).eF86N=
b-+dCA8K\QO1&?b6ed/;e<6#;QFd.M0POd7NM<4G[N@F,C;LO3gdKbHKGGG6K#4-
27eD,;/OFJaL3(-6b>b(T50-@M+1CXY)D@-fa4G<F(U3geZ?]/(a/D/V)a1.^2-L
AUgT;dNE<4YCO6_aafC#??a/^\_[d.VL7ZQTL)-Q&I>[DR,;;-#eH=C<d/K,#1XX
PM#3+@1f>&B)==59MWXK[F/-RH:EWHOR+)FN_&FdQc5IcK+S6eM;9-AI5<[08dUH
EFdZC(UP7JM<dS3NJOOT+:8[+Q?8Q5@f_.7O8)Y/ZN3@6(:[5W4YdCe+SI/\(0S-
MM?6>EI\7VNg>KC03P1RWK]>S\MUT[g+S3LJXC33ZEM&A7dZC;9a+-R?14L^+CKO
Ca2B<9?9f#)V:L2QM(RJ0/D/g^W,D@:PM#<]M78MIJD)Y:=cdPQ-UBa1_&P,0@^;
0?.N[Pg9Xe2QBQ)3?STRNVZ.UV.GG8fQUdX_,<8faLQ3ZD^D7>&F3+ZGUA,&/CUJ
I6(_]\B(.Q53;M<+YcW#QWW_Cab.K>RTP-DM(?-XH<gUVefbe&)/RHKFZg4TC)S#
47?M53OOIAE_Y0W:DVbfPP;Y:CAb0F]QOIM>85@Z[UICZ=LaI=2YfJ@4A-3UcQP[
L?cBLN-_SF]L,.@b#(+APX_3X@U,gWT6H#fZY/6WGHbb-3QMR&4,20,[=+9Q_CQ6
gD\(f?@_2YF(WH9N&+DS\3Wc\\6GK;8Z:Z(g/MAOBXP^_bEJf[@6ES/;-7S<OM<1
.MM-UT]e:Y_G^-1V0b@(GT?;c^ND(Y]Y;1XRZ1/>#<H^6EZ:c]JR?K(VdT8<d^\D
XP:.@XN_C;M@[#KD:VHQE.8^S2J.H3^Mc^9&;D^KG-/fR[&?28cED>AR--S-LZ.?
BUPYTCaYMbb5I7YZ[OXa45;I_VV)G?A=f[S&Q;8->dZUd#+,GZE-DY_3BGa@J(ZD
C.ICXL:_&75X6.UQ]d7@I_JeQ,c/E3/U6eb8XG.:REBPO<OFXCZc9Xc^Ca]/GX?<
_>&?(KAdfDB+P&=H7Y+&?<,,018;g#\X7YQ<=TWC^2L;Pe<_\#9VOf2=.c=?aO51
?9+HO3]G1<BRLD:P^dL\.PG/DcLg^U+&_0X/5ZEH-Bf)K1\Rcc2TQ2G7\HGJ9,;a
.4Y>BKNL,6-U-dEE/DdVYdaS.F/IPG,^Sb7g2Ycb135&,IH8QHF11-@MEcE,][P?
<X4[;eZS^deD_@:KL7V?D_FSP)GYGTR=?IP212HRF(PRd((I78@#C&LKPc7QD5g8
NJOUfY=_P_3aJ]\?E/WSBZ/)BDgFO(a0-ZE>M/2HT[/,]+cgCK()MAV1M3:,(D]/
_0DBS_;UI?c8:E<M;^4KfdX1,^gaHH]-H[+5(MFFRf&CBPe6Ob&Hb1<YZ:5)HWfU
MLJ/L>cRT9NPPVd#1.aJGI8H)-7]^I(-L3JR/3@LD@0LbT5ZGQ7,aNM]>=BXQ]NI
1M76H).N)=GU:/ZcgY0P)QIT52IW:(1=#[C0YMD.VY(>J0aaWD47Q_-a-G9[aM6K
&L_W8Fc8HQY4[I5)2d@>5c)O&?ed\)GEYPF(>Jc4>V&Tg>FQHG5_[E5\Y.K;]dgd
<a&f-,^EG19/9DZMI;FDZ(C.V3f[df7C9U\P/V]^WGD3,1K,BRG@(DMP<7BD3QW[
ZVBZ&MXMRWQG?Z<bQb/ZdCDIA/\0^Y.L]8\f,fL[@?OSM;+J<,X00G0UW0/+3EI8
Bb8=.8Xc\YO6_=>+8[VN[C<=DB;_^G7>(Gb@@U-d_[YF&aI+4VCeK:\HIISd>_O-
Y4@d08WZIZ/^9&Ie(b;[COV@5XPJD[\T7\eVU.L8;&Xf3(^32(6f@MO]YHc?,Ie5
gM&8=3#-6A60?N+/++#69ZO=X@;I;#cRI#YKG);&UF&Rg:W)QO7.a#U-9,?g[2Wc
d#;)F(FXCNF/CBI<Ed[+)b/G]dO>ROONL&Z6C#[VPYGaWLd)\d/IcIS]b0)?K[]C
I=N_,)K-JPbNC8I]GI\+HIW>;2[3G#M5A_3_P(?#(Q/5?G]LT.EJEF;=<1+NW(K<
8c+X..e#(E?UMcg1Y:cG4W[Pa9-?@f=W@^GGDP;SNU;96)8S>6W&c/Od/J_+2\7>
OP(>KJ)d9g.3QHCdEM\aNGI.Q)3LO3-PYBW]BVcO#NO;Q9_12R4?K;;)LQ)1R=P;
<#:6])Q02C;?_F<#VLD#3N.JX5=OP(8JPZJ0L<5Y=Q.0R&+M7:gQB<3:G1U4?.NT
-54-W&;8b,fLfX/WVRGEPC^,+McVFCV&X_UNM_G&+0DZG\/H9gR\KZ>P?Q02f(6E
7S+^R#Z_@f(4J(J,)?,DUU-AC9MWG[e&9f8CbVd4_ZG3^Nf5ZLRa..:,G5M#IKVV
-^D.aNQ>R6Naa[LG>G(@W[A8cMZ<-U/.FWVgL-+e6ENa]O/?;0&G[9#(6PI/_beY
MDY(YBeH5&A</7&B&Z[-^--?/LQL_9R24=3>9fH&b[)]+VGIX_f/\0c0\J<e&68a
613-+N)>d<,91YT?B(,HW@LX7V;LX\MMA9>dPS#@@N6)X_Y259:=:,T)0\YcAI<J
@HC/JU@QN/L12cQ\\+BME_)agN/#&2dYU=RQQ.\4Gbe865A\=M<3V0[^/3.gV#0)
IQfC1=4)A.H+F753XXfLFe6@D0T4Q,7BU-C)1S)5g470b^OAbLbf)Q3_3H/;0Zg5
3POQ40BA)OFe8f.CA(V,E0cTE.0=M[(ZC9b;74Q=#KQ.&1VW:.N</QNFAU54Gc_+
#aT8XUdCb4]ZTW,8X#6CeK8cKeD7H3:c:NMO^)WHf[TKLfM[aPEeOK#.3E@7=-K=
OeN[_P5TWDE&[?63YbZ1)M\OOe9+WYKHTO6[+TG^6]d,A6_U;UH4K[2#2)A]aYQ4
#dKC64XW-Z(c[&Oa[;TW6I,RF9PXJF2QQc,a+\d_fKV/IZK7B(VE0a4ID7&U:C:H
A3aJU4>[;YCbC;^.MBJ:,L?N08;3..CW;@d?HR6/W@.C.-f\Y]N,SOOJ=,H7CdZV
+<@(;5=V+T/5F8P&G[eYIQ76#@ZASVf<H_Ee(POIO(OUG.2ZEBR6YLe&;&&/31+4
Z(e+)N>PagW8AF]#J+6YbQY(E^Lb5:dU1b)<EcUCKf>8<#X(R<)<+/1EGWaWJ8Y]
&?+9b-W<,E;.?eE5QRMUO3=P2;T97BKK(dDf:e.F/KdM>\NNQF6.LbaX0JUVf-Gd
b6^EeRANZc?IK-#,c<KNI:M2-(-9Va)UW2?V^[YE^U9(FaHf(eF:@\D=cFW//F2M
9.>#&((8U,#DGOEE=+EOQOH[>MdAEW?+4R/CAdS4FVYPI78]>9,-AZ>MTbN#7X=3
/7ET;=(;6B:E5LG>&;UCC)>Z_D8<bK?_/+[X==XW\Q3INa-H\.V;K3U/BeL83fU5
/8=LH=LJ.IE]2XS8=8c)1(G(d?>AbM)aP@YgB<)Cfb-(Z#9P_Lg4D<&B&6V,M4O-
#GMgIFRELJH-GR,GXD0:cLg)MO843.\0d@-RYg(F&PU]L7CSP?#^VWGGO28+Q-2N
#CD@T^5<7#>:>;gT0?\d/N4/IWP+L6YTGSQ5-=0J9)&AS#_H\F5dIg&Y@RHL_=d0
38>[/W6H,XXINFabedTR>La^TdQB.QP/T7CF50<E5JJH0Q_^\WAZX)7Z\B9[/GPC
gD\EX4[3+>\+),XQ@5fg8cIe&ZZFECe^2<PR9YM<aB7BRG;:WD^eG+b4>;/;>P[8
B+,=++Mg>@@.5YNEceC:@A1e^:9\gb6-J;;;EIFYR+gfL&=YKZ3FME#]_b+65H4;
Ne63DX[V<&31&_>H4ND_?5-A=4&UJ@Te^+3Q?YN>)ROM5PQF+UAZV8K36[F-C6+2
G_/GS3C1fW_4Z@&^)F5C+4W1\4T7KU=OWa110CbYCXN\b)+M7S^2ZQ1ENWe8GMKM
@AQ@7MBXOgW>4VHB6Rc=\UfIcE<#Y^9_LG]42V5baU?RfVG+be3\a\Z^J&>7&)[:
D0\:8)SA5H\XPba4OSB:,dS(a>NHGV3A7PB^P+<b8M]?2JFVDF0PF&BEM]=H)VXU
NW&^TD/K&=WZ(PHZ@V<,QO3E?_O8BS,/)Z3F8QAXMKDU5M+KN^QBa)@@B>M_Vb.[
B_^c11d0,,-(WX.+V;AUDQG,?H;2fA8H4fG,B^Ad4eE>dI4eI>J++V2)&RORG^WF
dJ)AB&,<M\/BG;:0YK^5H)+0J-EDCT8T1#c,40X:d/43_A@ET:(AQY<JAHU\[/A3
].I)1]-c[/)R5#5MI82?L&2FP36B;#XC?#0T9Yc48Tg.D2SB97)2Ed-T1cI+U_:A
I;fGYMAWT+DQ?cPd\9&T0a;GDL4TSbNb3Ld,9A6Tc#4IHN1CBYbfV(,;2fc)J7=)
f7B[)R-F(RK2SR\a(=JObR=Qb\Ee.YT/D3:.CO/]\L0QP=71UKeI]Sb;^Y&cV.=[
6eM0DeS6C(;+AWOg?^<RI4.F0:d7RF<=dF:4_TSSQ_3d^NJ^Gcfc^LPRN/\B9N>]
A0YTN3Y0CXCV)4]f_LdB@+P;4gX6@A<<_&^MP:ZLA1W8d=[Q95AI2.g2(#18NBO4
7Y&VGAdg/AGaP1d3b<W#Y2aI+&DNb@d;<@_>A[>H]+5+b;Z.DOX)]bd30W97fTP@
KeGKSQfc:<^e:K7Jc/Y\DQ@S))OAe6R<<66&O8BUZa<3fM59O2U:W1HJedA5)M/8
0?SU2.O?J8f&b7eW-b9DNK0eOf?>(@6#d\a#DM?94QgK\f\B-]EMg+@6,\),:A@F
6[#Q4:]]\CDM<17KQ[<&9e1gN2&YaT@2Lb;V\VI)dBKceBGJ6S?&Ue5aK,R:7&d]
RecSb]0QfM52Z@+,L5Y@;?LXe3(^&7GPNcB:HW)WSNKg;IUba]/f((\18W4/c8PW
UMB,/1Rb&]?)XW\JX5TQ=/B0J07J)LYWbCWgJN=@\&L/.g/4G@Z/IbRV;a1A9R)L
B_JK?Gf71F3>J+=YK7^7.O(9ALONb^@4)-8)_XY(8=IZ;XdY=4:@g0U\9W937=BP
OZgS83J<2ZNNCZ1&d&4>TEHQS^2Pb<LLAJ4:CabCZGAgV(cBE_>=VSB]2;T?B1/O
AN>AR6P&1YH1>TfJRX8e<HVZcS6Z5cR9OTJ;#B/FNe^AVcP&=H2F@[@870^MKWXB
C@&;8U[V;>GK(:S/TAgQ_@<U)Z^A1#5+YOXGU@fE=M.6##,FZ87-TeVN7]I39]LG
2>VJ97>[I?PYUPG6?:1I>/2OT.T@T[3#U.K[(GCOQDZ3+A[X^4FTP9Ge;IY_EX;E
gN#Y>e+Ob(;/ePSeMJNE5880TR(X5K1JE7KO7He3TH)95KbDMI>_)VLV[=AH;M]C
eH;#UGGM9?GBS+?)[3>RX)@HYTG0=.e/^3b.)@A(8I_KFZ:QEHD-M[\97^\2U14#
]72QVbH(JC,JHSd)S9[M^D0cI3/3b(^U=\e-MR<\7f-?69<^V_5Td_QOee+PC6S4
;+?()SED]3KC79HEG>AY=]]eWa.OEY/NXPEQg<g(7;eQfR)5G+Y@-dNKV2\E&Y5e
b8;1;1=MSME41V,><6L/^LO@7Cf8e5A>4[]ZfeV#7<2;@b]<2/g>EC0CLFVBaQ@,
^U5f\LY?^X2ZgRG#@)EOKT)>A<ZV<fX6a250=P&6WK5L13770YdVPe4&]-#fN,Sb
DgQgEAZN8MW?009RXFY2ZOZE&_-W_SXC39-T]F(E.2;YGA(Y&AHB?W;-YCYUYdJc
eU_GZIF)bD+-0L.g(HWI&91=_)1dXg;:J<HRW9-\:JQJ,AR[F[Pc_8<Q3fe&Hb#W
IBdI^=5FK.B^@YYP,0e8<J?+1+@WDeY^fFNfI1e/dE83Y0b4Q?VZ4_4:=VeF<7[0
3.51D4^>[0.?956>/1J5F[OccGaB:M:9]2O.WfC&+V1OfX37&,cdE<<?-9/87^9g
PdDM?5IOG[VE2W0Ic+QP6AG9V^:7H:aCPB&I,+eP]XY7(G14:QCT_X+[3geKCN1G
\5]c_[?7JQ[EaL+HUH7g1.6]e-L4<^.RZQ4A<4^0PI]=K^e=I@CX_U_+9Q_7:P.(
NO>3&b3&[2N/:[^a4ZR:X0R_LX8;BbXZ&f7@/MZAUA3E7E]b)=\L\KY<^<\H:dT6
(Ncd[<)Y]8<0=f0)_b30Q;4?O[IJ/g=O8>02;PQSd9]E_I:eTE.;fN)TcU)ALAX&
V@ac\/aD@a2FKL^V,+&ET27K>bd?G1&CQegPWb262dUGA;I<dW)<H#?<H^U5gHDD
a4,dFdT:EJLHfNGG2e7]0)HZGJWRC28@[5YGJA=,D&g?dCVVEMK+-GRfd&7P)1.;
\7<(ObO1g#f,8WV59=85GH6NfXELg2;-M?Z>?3AbA\d@JHa_(>IJ:VbBC(b4+bN1
dJT,UK-.S.e6L55?Q99ZJZX5BEK-ADT[<U29LF8ZEbcgO(N46_Od8aL8d^M^<--4
JQ/N4Q<L:8:AXH;J:PaaW-J:7;B>X;YC\._C-M^=C\ebK9&cHQIM);#aRXcC>aE<
?1\dTY&aBaE/39HBMBS,+EWWTSg-K&J#9:3ZE@DF2LDFOSVSKe9<G^.YT<D6Y=/d
+=S@MU]S<1Fc-dC?<#9_=LLPIX,LR/VHa(=LePGONPK647d8AQ[Z&59#DYBZ\BK0
C31.R=fKAX0A&/#.-a7(=f_9[MRa3K>T#=7-bN9,F]B(Gb^DW_-/48>b^5^N(O_.
WV;=4O&I1a1G1ICK]a\W8aEDd^Hd,MZ[g19.g\(W?5O34\OeA;egJPc[],8?=@92
]d[SG&MB7bA]4e04RX0V3@F953WS2&=S;HE)WQUR(f,@F51aY.G&LcEH\TWW<>7^
.O2#Z+3[OFA#Rg8C]9@K2\5^Z8]WE29gTK5ZAVG?,/#e4S>_XMe>0D-\O;H(C:,e
F(/&bGW/gdZ2PI=&0@+7^e##Q(A9GIUe+/gC+:3Z0@3#+V]b4W3,)E;N=I(5IGEM
,LMe&QeM?ecK4Kb>@7+PQS83&>E5aL-gAWYR_Xcb\;(X.5#QI02?#.3AW(DbM[Jb
c-[UL:=VQJdR<VHNCS)VES)C2-082<##.6&GcCQeda3-(B8B[&.c:[^9eZ;IgN(6
cd18cPBH(+0=#>YA)UA8c_K=XU0]&Y_K]_eH3TGa7JZ>^ZX[[TcM_@NA:6a6d?_V
A[>9#MNdOc1]JJCedH[RD+<AE,9>ZeKQ3/]EfMH<3gUL0^N:DacD;COa#P8+9B_=
M5POL#2L::NFc3F&IN@)XGF@aeQGQ]>\CXJ54=/?\HfcCdc@39Sa]TGW-7=JXT)J
+R@LV:7_/&Dc[Mf#2,M]SE6DO<(0;?_Of->VKa15).R.5<gFUD0-:](NSL/Tg6g,
?WPPL7JT^D78>I@&^\0OcCK[]OSFeVHNG>:1WIFU>OYW>,g-;)JbLLg:.c<.+_0]
)BVHVNJ4CTK8ZI0]F0(NHYY++.?Wd_&-E&RQf(ARc(5^7EfEEX&E^PMK&O:#ZL6Q
7W8)XWGP&;DfT0K&G26P2a[,W5W>^0b.-#aA0#/NGDR6>DF#e:dcdQ<N^^,Qf+,K
a3T?;B&aLRMa@A_AYS4)9gM@Y]0/-1c8)2-&;SS1ZCe;8fCc\gJ#Y8T,5YESF^]f
PTc^P)T+eDeF@O>>,dS0E79d>&>;T8[++VL:CDaJ(1\4W<_=Q.M#gB<He[;L9#T)
8E1/;>,/07-g=ZO[]K9R,OgOD^;FR<&c6dTNU8g)MHc+2&TdG</I<24IG1<DL@[R
A9@e.Zdb=##T<A..ec)cT\FfY6=B/=dfY]1\-U,0/)fC>Z?KDNHFFc(R\Lg9bJ-9
)\C70X=85GBQ,=Ke.,IFAANfMD[-732-aZ^bV:H:_(ZZM)eE0OT<Z?K6PLB?-KLa
NKWI6&e5Z=.a=@X3;M;UXEaT,9,:N@>,=7I[/C=T44d&;8N&Z>;]GW&G-BKS,6aa
I<>4#_);VH??+LE^,1,YfDSGfHIHY.d[0X\VMdg#XX8Jb&]FJ8@F\RB/a@BgXQ.6
OMHO\<R?g.5/91HgO\DPV@A@6_<KZ_AY)D#;gbO:P77O;7>32C?YZ)+@TJ/T])=O
56cfb0N/A)b-<RgT&f[B/c-]_Ze6eLP05PEB8)MMcd?GN&d<]=\P.@C>.1a_OW8M
(e(9\MNENHIdAVag\#MQT/)N@MQ<a6V30.9>I8;E>NQaVN1Rb[I=a4F-aSG>334^
J@=T0=6R,70bHIQPC>aQ6EV-D2^?>]NI^Rf1+8L0P9gc)3U&&43J1c:5)cgLAG0^
1UIA,O0PEg\)702\NM-T1>WHN?GY2:8NQ_]V9Q2)CJJ5S[Y@UE[e?HT^cX7:d5W;
V4?UXM@-\;]1CL[+HAbd@<A/9WLU3-K.(/gd_O8:=FL@.?4g)TN6JCE^97c>8=(8
g6ZZ7]DW&MQ>g^)8QfNHVEd+.,3HB2M,&YT\BQ#VC@?BYQHW7A(c;5.9K7&P0bC0
-;V7KIL6<\EEf[?-J;/:=@9-:M0JeaK&.-1:),6A4)eUJS:K[\<cZK?6<7CaAF:R
W,P#S8.7Z3(P4b3US(FT[2^?X1OUZ&:[+&;0E@DU_+-dPbT.d/g(=gW+BQ85Y:><
6L)Hb\Ab^Tb)AK;4gO00,g1\[eDgYJ0MT_K?CCK.SW0e/-9IVG)C(fFPVQ)3H\If
]ge@NJC[/W:N&DZ.0^1f]<LYS&B^+b7^8-#Oc-Y>]1Sa3e-@GK6[,?OeHX).NHgN
;Y2AMS>M#Z<BAD-b34QJOBgY-#N6FK294NC#;1SA4GDYC?;(5:KV8QKT20;&F71<
eb(]72?I:Da@40bEFB(<gNWA];N5P_aLM78C&eSFX0<:L3/U:9T3<dU+8O=T1_-F
cM;FW-/N=7WLGbYDUY9I:,(PbJaANIY1c^K7]\[@P)RCM8MB_4^XKcFD&2W=fK_-
.6_,FgP>Nc^?R31OQ]I1C[6gZ5+B&5Vf><LLa=:PN7_LT<1PY9He95;:1aRPbD-Y
[1H1>&>)M[QZ-7cU9/#/X74EY?9>8>5-7W2B<)4GJ+g);^+MG;\AY(QbYe]IK<-+
7Y3#<__agY3e42&=H1&YdYJ/T?&I4)8GJYL3.>C,@B=]B@>F6UFcC-ENBR2[71?K
QEJf4EM#3FeAc=2Jf^_O7gBd<@340,=LXZVQbZ\1DN?O8H_?7AfED_f;5A(Eb9T@
TX&.]KbKE-DObP]K<]JEg1;eX1E[UEX_Y#OY]C@V0d@GSJf)T4HI9<(N__UNC3RM
446I9]/DZ+:L.3LYRZOWUOTSeZ_GF9TL_WUJ<A)Ab6Ef.Ja3&?>G2e-<;T::2@?W
__3>-1I5X/4[\VB;+FB9_S>ZC8Y/=#JR&;Pa14_J<.(7V5aKY2-V2ZRd3I-.<ATV
DcNS@26c7[]Ea,M1NdL)K@NOA2<BaG./\?5HCgF4OSCSAI(MNV92@J_)7076L/>K
0?135KA@YPeFWRBeK.9D@^I0<9d\FV7Nb8JOU?]LG_S??D5bM3,V0V\KPR.B/=6c
d<SgR2Y)g+=91;.g(:Ze#9D:Fe/3P5KL=RXK]_-ZSMYTeLG#[9R=b\#IF_U@C4(K
2F=<aE/4T[@cWe@\_4JWb?HRDM^0ZRIBQ5)bG.MZZG,_V:)W0(?DfKcP3X]a79./
;bXY83[;eJYHT_#O-b9._g2?/:XGDFZ52:.1eOITGGdNTE:4J\0?g3OLIAW;-68E
e1I@L,=Ua,FL/TeC@H_TNg/d49TH4T8&dL\9SEXe&B/-:d,NZ5LGF9fI4cYf]&0(
>WDBe@-/<-^P[OUG2,+KaG:8fXNMONP>>;6LO3:(?Z;N^90(X(^1>-aC#R/9?W]c
S[9(L(@aU61Z2Q8]9&fc(:/K93NGVO7?gL?[>](6(G/6ENXe(cM^YIJD\gH\1G3?
4TPKEa[9-UHe0M/_(J<&Na=D8_>fd4Z]=3(Y[A6Ng?Ge1:5dG1f^Yb9+Q[eLeUH(
8W<W9JGQ5,40cNeL6#X=G_gB/O[UK9.T[?T5:]IZR+35P5fJcda,#7Q/ST0=d7d>
&KN,0Z2=AU9JPN@?JWbeK0_WHcI]LQW.\_;X[XC<8;=Ag?(\KVIeKf0,YU@[B\;E
dQ7cS\I;3-R^C=;BY_S&.)66S5_S9K_KQ.6Hf]HFf<A4@/O^ccd,6I]0RM&[5HS0
ed_Z>QP+aH4;00S=5,NPZS?@c2+<?=Q6Tf=1,ca^H8Z&.\U)KV)aM.H)=&PCSG3B
JI5)NM4^JN.6G:5V+RB4G4d6:@HY6#4/0/aM4-4]:b^?bfP?WVK23Y;UCdU/Bb0=
=eJ<bZ\MXaFKOF1fLb?OLKP9KI-7a;DcSRC61Mb7R&7.IMI(d=:_RaS5@d^)4US>
fJWWNg[?g;G^V>B=XY0X:#NRM7?GJ-Vg)NEJ2\Jg:Z_aRR2P@8(CAHFJ,T3O33HR
)GC>PFe<_4?[F=A2G^PPFOH]]NX1bDBEN,TWW,YVNHb6\^15GP5U.Td:11HO\43E
[W4b.>\\Jbf7>HIS7.;K15[HYW+S6dg\/eO>L,RKO\:_E^5&4U:1Q0f9/:+]b<-Z
GYPZIMU4^O=C;U+8<VNJONKD6SfX3+JIG_J+b3a=@CC7S[Y1J^=^TBMPLO3K-_1-
_P)EA=X/:>_edYP[^@&L56SQJ98c++T-e\>A(J4BRbZ)e^R[Cb^:A;DN@+HZ5<):
Uda]9J->\KOU8V3,P;:FLAI>8ba()B)J1AaU/V+,cJ+1?\]VEfEg5\:WNeMM<>C.
D7fg,f&#EV,GRdEBPJ[]B7&A_;AHY4Mc,O.#6U(F]]#=2?=#J.<3EXX-=.,G5LgB
<@4a6UX,)Pc\OJ5Jc^)>?2bdLa/f&Y5ddKf&XCZ>_/feTQ[4FEL:f:S.F7Q/24+0
_Gb^>1(2+U#OINO8?++.Rc4:@2JEZV/,>PZ,O16aN.,ZVLOH95YYA+H\J<cK_cP\
FVP3dQJC-D8g>Se<Eg/X[]Wg)bNE0MW8GB9]-KL=<W;^=HP:f(]6eVC=)#/&+1QC
#5aX1\2eQVT3()<OPB+@>MR6e<3]:E])7-U;1K#0#9R7EN=VJC9)BEJGD5c#@]Rf
7a?.D6T\bE#39&3)9>HE[0&aM,553JbUg)B:G1YEO]6>E>Z3];:P)I-^K?5WHaAV
/,Vfge8O\Pc]ZC?aRV7HBE3/eW2E_:HNY<K-55?de.)PRN_]BXA@.N8AMC@25QD/
c5JXUYaW-ZfdJAc;G>RdCNL>B-+S[>V[FDY^D^.>V><UY&FNcSA@0^[ZW<2LF8ff
H)S8g+F4P4DUTDH&@M+:3RGe\I[[)9B]D1R(7Ld:,VUA_A187@<,a&])BF;/E6AK
Nac#AV7eB3NCa>Yb]QPG,5fd=G(gNf:W@4SJN(d#0,eEVNZH<>XD[SW8c4:W/LZ,
dFHNCD+:P:CER)BA#EN\S^XYAW\.LA7756ZE<R@WFef[9G?(ga1b;Y(]#cPNF_K=
F<E9gD_dK7#a>TDe(?+T388F4fA7/_>C>V^e/L7DM4c@M[Se<-,4b=MTP#?B/J?O
C-DI<F=/W[Y3M8JOH#.g=>d.BXKgABL;Y-HC&4eX268bD?e&L[:=WcN&RU#T8d=0
PY82L(6O8+[A5>e2CZFBbJN[(BC86A-,5F92M]=925P8/5MHZ:a9].1P9_b2U[3d
=I@f6AKXdR&PK3]Y\S3<a,3>N8Y;+1(I8,8fS5X]39,;[IN+YTH0F#4DUQC->9H2
OUf^9&Ma,6)64,KYCaO8#]/5cV20GS;c924\IAB\.>:Y8LLX9a1<LG[:/JKP-WVU
#C&T=@NP)0U2bBd<N?f=2@Wg6@0@U_5,IK71R1&P6KZO68:\B:^H;]?6]4T(8XM&
Y/U@6?IfAKgVA?@D@K6SP#]b@8^&RY[Fce<PK9OaTR+&G6.N)5g0-=E/TFfe35_-
]NP20Z6C,;W)c9@?W#1ST/eN;bHIDY93gLeN6;@G#WJH&QFJFAKKdP.#I]8,_-XW
03:HN:QXGO<+/_+EUQXRRKNK<(Y797U2dg>[0JE@@N-8&c&(A1g8-ZCf_:L19_[<
?#@/eL#cSfE0M?[bU_49a6#1LAY?/P:9\9+#U#gaDDdZ2c64[I;#9LCW55K7TdcK
YX=ZPRTOeO4P\,fBF.MS8ACb438,g@@AT#L?He1gBUOgK\N;TBgA^e@SRHdg(5&@
cI.>T?a()N.adg?aP6RP.)T:;[2MRHB2G;5>1HW@QAXZ2)F9e+ea8dV6#V0PD+1Z
3&e+L>Rgf]OP[T,FS#^-e^#7^S@0YHEg.\5H;edIbfe4#2?&=QVbP<g7&VY6=S_)
6HJ>>a&_cJ&-D3>8D-RO/8M5R5.WIW+,?TUI+)7T#\Bf33^PgdZR;?&323GQITe.
M>6U+P(1,+BH6JT8&PcGUP(SHMAI8&W@9JRD:SW#0?VU[C^6^Y6Y]6(91g7.gA>&
A9Z,#;F7-^WD?C[F];JL42]#aaRZ7DRJ>@>9+1fJ;Z(a;+6(/;Ac0<=>bKI-EPVX
:K<B.ZZE04RE.)]bBeF26f,/8OAe/XREM1Y7X@N>6E/^.3dG]N&9BGZa/,O;2ND<
47;<_TCD?E5[X7d2)AC\:QeP\D_63G,<C7b_#_Re9RI_eFG_8Y\[_BLfgd>W[PYb
e8ZF6:1Ua.JFg-O)WZR(C20,Vg]b5HP+&QW+L=K&P[gb)ZF?@B#eQ;E)9:4E]MWc
7<8RM[#G#U,T[?6b#S?4?A6AP/,f>5?CU.<+JdQe]&(Ua-f_JcUQ,>HA.#N3RPUf
0H)SSXU5?G&b2#41,4O5[&cYe8VO(3ZfM+=,@?//Ac5.5-&1K&:2]791-d^HN\^I
.))>0A<Z_6\[/[2g^9<;+a/^g?0MKU6\1&G-2WWN4X8FZ^[YVcB)/]XB[(S(+dA-
?28Q]G(1Z-/VfCGM7_RJ1F1d<2.W^H21GZKK/9aF^;C_M759:\T2N5@L5IHA2X6M
FFML57[7ScP1Vc>N;73DAE&&2dL#T8^70HV9>UQZHH0#:,S/]=b:b@(g?-VaYgUK
_C)G.0DgcC5eF?I;?+7MQXA\,[IX@>K]28bA<+,SC@AHPKNS?Y_Xg0ZAM+b,Z)8S
\\,46NBa(N=d?JY]-IV1?f1S\UWQ1:9-a_.?g118=7GXMR>1fXOVGf[MY[Q&[UR=
U+B:J-eOH?]JN[)HWRE)IJ=SKK9b@7<_/,V)YO@WYP6Uc=D)8WQ\]^50TgY[]O]Q
24&V-F,,P,c0\90#,/eR.T9K?[LH)X_cbPVSd2@UJNHfa?7ReA2(\2)IL9F=LE]H
V/YGJ2Y]BA<CDG3(8\H]_I?^E:OSKI=f9^RTc<cS=c):Q(&B,QWWZ5?<.6N_3W\J
3EOM#DIKC].-3QHR8UX\]VCJ1IHFVWVgUX@S&G7+&Z++@9.>(A9?K2C7=G9WS+I:
,.1#>[++d<B.\aaIUH-N>N8V@Z?K2TC,CaX\A.1.Wc4)O7XdX+MFOYBF-V99+/TA
Ad,3=OD/gUTRg;^].9A.D;#Z;YaV)G^0<E&ed\93cO-Q2>TY(VJ63g4e^ZT9?>eH
V_W8^[6#P0.a#99<1PEI1ff:M:&g422.L#aBCXd_S<JPA(\O.Cab7dPAK0GQb,C\
R4V>;>:G?L69fG,0daPcY9PX_BA#E;Lb(+_#-FY-=8[aZ.:7B5G.@<TGGI#00S1>
RSMG76fc1IVK:DLTaPS1.Qbaa^(d8=+_@?\;dM4-@&<.?2>[8:,aQ9ZBA+^3Y&g1
JM4Y)W#>/-;6]RU-2[I\Q[@AFE83WEe6012G0)FL512#WMa+b[YTg^FNE\\9,_[a
c=d1XL0,d/a3@-N/ZfG(VbS83REaZGNe?dTa-BPMg6a[(-3C]gJf6Y]7c3O0RB/P
>aIW\SXT+Cb^<c^J+7KfdJ>eG2X7H?7&WC:^M?bCK]&8F,JZ@MdLO8@69[BYW)Me
S5f9E9<-A3QFC^.D[c.F4g)-?^V9<(&TJaQ^WAbROS]3-<4REGL<OF)V?7G/W9-e
,9I_MDbgA=7+8X.W7(^M\a)fUc7LSGc)Y4+:N[aOTDFKB_TL<)\NB2&0P+Id_B<L
<U7XJ_:T@+<1f,IHcI_^d<T4+WdFM2)Db.W+eEMe[@EAD5.d5HCf4?FcJ5Z_N3\L
a>5eIa=ZecXYEgN(\0<RZE\P.8U@W/d/g5:W(^G7((EP/]g;&O3Vb<bd^@A(N@J4
R1=I+[fYK[>V<LgDQe.c[(fedI(STe5VBbMF32W:]E[&)@MVW6gL2[95P9;4-ZWD
S6g,?0b=OdK9-;+YKK632RXN;0P5>J9ZYAJAD:7Pe6Y&38YS[0#f(3<3.R_,7\Oa
Of2=T@DXeO6bD8HW(O:++00J8N:^_D8V<G9VNND\ZA\a:-^4I.bI<F<&+9,(fJdF
ZL\0@-Ba/53)f5-DS&HI@376YaOVf+C]U0/S1Z.aEHBLADCGUSaNA\bSB6T6-F,(
MQ,]HHT]=MSec.L60<1gKdVU^Q>3d/Ue5;A;0B=f7IE&[#E(->cOP,6G+Y_b^dOQ
[a<>G\GZ,@^X?W</egN[NQaWYd^7ZY(-)R4?g)(eK6TQW_M?8.W#?U&<RfCJ=056
-gH-T-Ig@#+O>S=X7fR?CgUEg^YR0Q#E#JW36gW1C,6X-:@Jb^0W&)O(>gFR?7R?
bCPJ#Z#Jc6\?&7JW)-MGPfA4T<?W:;D7DI4U?fMHL0.Z0GbDaIUGY&<&cI[1Q,QT
7H<79HT7K>7XE&3g.bXDTGG70H4DTe@F+c42.[PS&ZCPVbD7C-FXMfP;[<-)A\8V
IG#U0XS#eY=c;F-V^&N0#RcGLFPX1CBb7C^Z&Z=:TSOAa=BB0=<eZYF7N);#0QC-
VJbFFL/U_OgddE?J)cK1HOQ7IEZ&[@^:+-/M:D);/-N/&^9@f3gggeDOQ\=32QIH
,W2Y<>Q<&TFcJD_(BK<C5H\P,Va4TDGGL&aFW_3S=e/aSC;((IeB=^ZV2B\Y6W(L
(?cFTf[bW[fR7c1La3[QWIPJe1L\3#30T#JQ([2T85gS<=&U#Q6_L9\P:(B_YcLd
(C)ETE<R7+Gf57R8Y2VFXNEY\9XG\5@JMIL]V1IX9+aU6?H/Mf;#>9g&dAL-UQfX
=TT_3g=VN]#]N?P,fM...3?G6X@);eHHWK3W;cf_@#U4S(fCdSE\1]I05W4c=1f[
./g\T64P)LR)S-^RSF(E#BY^:UF@1I@/TI0=/1dX)MOM+U)Jf87[M8AJ/HRYLLe^
0^D#S(-5bHMB-eL8,d\)NXUM2a/gc<cX7bA/3^d8HD2W,G^VDX/R+;fH,)OW>V9<
J-E(Uc&N8ag5[T<W:).O9.aG]O7Qe]cJ<?K4g>3da.O5RMTW(>W1W1e2=LF#2:8N
-E(WZ9XTZUPV99,^_]:^YTbT&bE=;,6O2NY;X;I1>ZIfU]-:IZ/Re\ZG61gGb0P.
&J[SS=cJ)V5A#VB[C#=J^_NRcVX+]KC)O3QSCUY[&U([-]GRJd]4(MePYP[FSEQO
CB.G6.RH6VEPa=8D4VI811\GZ+Vdg@)8P#]\a3f@_ZTJP6BB=FCc;bfJ_8K@K-5g
bSAN0=e79b;FB>=];J_/Q^)OX/B(U&=C>fGG@?H4,_F2(d7b5&I/8I)>53]RZ=^F
g4XNS[.0:15G21QLLENP0ag501@<^a#IY3_9E[(c19U]^YT&JMB5_;b5^aR][LA]
.Y7f;-SM=6<(@:dN5W)<fOUdIREXge-N?b/O#C=AL(e_fFY50g<dgQM2BD#6G44-
6/KW^c8JVV-.VHC#&KC&U_Y0KF34CD\=^8aPEg^0gTaa8N#5Pb79/]S5f.dD^UVH
UbPHfTe>XZ0=+>@@5)/\_+W3K&1=9[90_P&(Q^f:[SZ5[PA2E698\/8WR1KSIU&d
-@)A-0.3<NS1\YW)FI&AR;:/0YYZa&MPFUIW,^:eP#=:VID/@\cUIC+UYfSCE(,U
8a7Y+@@JJH\\A6L?I=#<bcgIVQ9:8;)E^2ecbd]SCRWJ.VD_9(T:[W<W01P&ZV\=
GPeVMZ<:ZQ9@YNP66_R5P,K>#K383&5H>VT1LM4-Q=LVK#YTQ=_aUHS0<WG5HAIZ
,GX0>QOF(0NV45D(.T(0@FWOe=;e,U-QPe?LeH]?]N:g3C]?CN?dI6b5e5:SBdS>
00aP-gMOaTEf[6M2/eCL3AeL11,M4GR)=X7@L,8]-[G_?OKL?&g7]V_&VGYg)#>H
9VM^596eUYcU<ORV@9>d[NF];=0@0DZHRWeN4ef=F1<E(f3VSF];<F][ag(;=4+O
]>JW(#=V:1O>/&G,UBDb__)?AH7\G:Q9\YGBL.fIH6T6>-Ha9HK1X)MN[F>V\I99
4>U>3\0>3Z4:O.C0ADe0#cOb-G3CcW&Nf.23NP,VA;^8+^#5I.a-g?15N0_3DgbP
QYWI:FYBQ3YdV>a5/g?Z\cO#6AaAg#bO#U1:JYU-QE,0#MV>H9W-/&9XOb2H/69Z
PPcYXMB@)IYD/VV^.LVDX1&aLG\B?]@^VV8-I378V/:eAWJ9&8I87RVH[V/C9^83
/10D5:FHWW.P/ZAUgLTDfb\BMOSLD(<<X^aPKQP=MAVUBfO#F1b=HY]6LR6,MC,a
GVZY:W1A5d\8,a4[\XH1BER82eE4D6d;OZ+;G+c-M5:.Y6TR9PA\VTbYP1cQ\@<R
9D-@VIGL)Eb498-ZKLX=KVNQe,E(<dfZJN(9ec]H+Y)\)^.RWL,L)JDd01G^0<f1
/=SO)&f)J\]7W+d/KNFX<7YcY)Dd\EM[]<L0F(DMSgb[g:(A9&N92TW:R>7KQW-(
Dd59^6dG6D/5]HPQO.e@?6c82]Sb&?-8#ZJGH4.BVd,^WP^C]:-gg@8,4^MB7#Z^
L&BBP1.3@BHDYMWY&)_:GW##4<8<0-65XIgYU[,4=&+44[E9;IW3YPE#6af=+.XL
aeOLJWD9.6GP;207D90+0X>QA6PG,M)g,]_N?MfFT5BI&bWEPNb3F3\9^-F]N;Za
-EM2=?LOKWT:K4ZAb[/N#^H7@9ZJfYMH/5R0T;\I9DH=X&)Z:@DICVJ&:e_,^_Bb
TFRHC6_6(RE^SO0HD(TMPLN_4/^VT(/JPS)-FHFTQ7E/:^c#9I4S#SS:?9&aG1Y@
XFL^#4f\f8e^<:WP-+\NVScWK,4,FNW9e.+?4g18M-3ON()Ra-8[#abRYN[9<<\M
X51X;M8][^MSCX1.5_B\e&;G^37eW=H/CB&f\4;VGM646g(g&#GaA-)L93Z00d4R
ObbfFMMWA)P4g>Q_W,#B_TE9U)_T_85)\?c/Y:[420a<NR\H#g?b->ZS[P?c7dd2
N3[dCR5_V#5]7JI3^FY?9&@KcV&Q1E&6WgceVK;#/?X.1=RCST4_8Kg\eY;Y01M/
>W6[5=\a8?6c24J]88-B1PP@C<UO07X8MdGE0VE;@]+#J#VINg95SRVcQ;M/3=H+
B?E-=G/dE]LQ>IdA-eG?aE0J;eZIZ:.CZUL)G/V3P;fX8aT0;d40Ba&(@_,^LG-F
R#>-J<:7592fKN;PXacCKOBU6J\G4HBCeQd(=X[(Fb:@Q=.[O0LRUF?MX,SY4\J(
-V38ZAC)/V(R1OCW0TD/?GAU[BQ83,a;Q[#OGZEdHSGT+&?dC])H1S7,;W0R\;3F
+@8]Y>.[)1M,+:@1/&K0d-3O9YX_;XW1_]@IT7U:6UKBdE2B??BNO.C/c<Z#/QCJ
&Y[N:61EQDZLGVe&9:g=OBg7P-W=WEA_O@&,a1QN[B=-8eV.J_.\PYWcLLSG&9VF
8FC=(3,^O=AINW],7b<W]BO:6MNA155JGG&M52HY<49IT),>f;QV<TX22BIfZ9K0
JR;=g/bVCNJ>0(32=?gbX9/#-0.]J_<18/\8b1FMM&4?Bab,a^=1Y1e^g<@V-Y-O
.-bAJe]G-P^cK_H:L91/XW,AAPC+4K(Y9R8YNX1?6>F#O@^<B,Z<&;a[XBOT9=U(
BR4C]^+#M+2+G3fAEJ^gLX-ENA>)ZO\)TC7;,ICEFL137K\TJPKdT5E;P:7.<BV)
/[_[gF&-+8bX@9<SZ2(ZUGEBaRMI6VcN.7Q4F4)<c:J0UQD?A]PQe3EGE5Z=bI13
QM_NSe(gV9I]H[DJ.MCQ5J;Jf86@?7?S/KY2E:WV9)&Jb,/Y,R0F)Lc99XHL72GQ
V3TPT.H3@JF(85LJNe5M]8:[9T?TBYBNZQ9W[XO?9JT,RT=c():]_=#71[E(+Td5
ac=6/9:2&\#1_TfYBGP:I\I2A5.33dA,aaC<#YT\=BeO[_YL<RG\g)@4fd=WdN8T
K@96#YbUS\U5<cE7,,(IgMUFH9-F?C@AK)fJA=)B5@R1Z@Q]O+2+g7-@S5P6RLUB
cU6FIO,47]PN8X7UIT#<@fXBQIfgN77QLJeK5UYZ;P,+N4S.6-A2IET39X\@)We=
(A/:Qd8.;&I)W.dPKSB\fD=6P;#_U[D[4eI(JZUNgecXYf;V]NIV<CS1Ia3-JJS#
2#EIMP]LPM7U_T/4DO(Ue.SfG&a9:]CH[61X^Q^.,0+SW0&P6.FK(.SR3b:#=AD<
ZNEX9KPKFgNUX.63[HB+2_+bSO+#+efADFcMQ@;e8[KcU2#VI+9V9DFX8V[RM\-K
^07T^O&A^9MI+<;1YLa=?b8Y>?fEL\(5QL5+#HVZFc3/\TX:/ecdAP^<F-3-f[0S
(<HC:\0dO6#2AZ[W@,=_DgMSd].AHMPLVgS.7Db5ZC.V2-DS.,/;&D1cQ?eUeWWJ
N(QI7N^AAHO,1@-JbJZf+M6+WWZ^)3>M[TE&<XKH23M/QL+_M_L8?AffK9+3H)<(
c_@P#2N9@P[3TFa5Q@QCe>HW:(ZdfP\4+:/Pd-9DRAR)_VO.79g]0/WffM6YR7]+
Xf,K2TOA\<BgYIA1X5e&=&R_?E3b2]f[(N2XSRE0;CeCIYE3A,^SK[CKBeT)Y#O-
bEa=XYMF,I>>8:SCW@Y)I:+f-g8&Gg?@T-[HT75U#YdEW>O0bbUEF56<CE=S\gJS
72;)a3@<,[@ZTNf+/XW&#7TG._X\OXa=2]<X809b;J,Bc]&TMXDe9)C+7^?E,ES&
0V7K+TVQ>D,IOb#aFC:^&_SVYSYR5VJV2a?Z@_,YBJJ5>?=&+Xb?6\f)1RGITTO=
K]QW_V23E61CQa=7:3N?Z&3I(Q_47AFN_RQ/-^IK1&41+?:dBf)1DFXQI]&RR&g:
(,#=U5()U]2N]@;6\Bed/5[4:OeLEI#=DKB1g(c>(#_01F3C.S,HLdT,aB/e:e]R
ZE\FP>08H>?]E+79IUN254abG^8C&R-92(T1H]&VG.Ha4644,668#gf]I2O@K1EJ
/_S;](X[&cM3_0aCTNZbRG8RRKZgHQG8CdebW8;+&O+Sb43DeOP.IMdO83VgT+PM
@a-DBETPLf7R2N:,]bFEA8FC[1_NT]=Lfd9/++2cE)YM#)+FN>-]M@/1Q8cYZ?X)
NK8<&B7ReN:FAK7eaE>\H7FSID:<KZ<VWROPHCa@EMdc;DCQ>47J.LP+3fb<)5c:
@/\L+)M\?YP-RM7E#Jf<dQAMZ=+Hg9<g8QcDC8[CGA=M-afN]O]ABOD/K\S\.^IQ
A38e@+&09T2-^5+0,9dXfa07aSAd76W7cM=P,4c-U;UeR]d-L8P)J)d(7^Y05&5d
PAMZd0\MfD^;TW\Kc2X,>L0?H7ZDb[XT(Y-]P@e6JU#4WGJ(F<##5aVF+.YJI1WF
SLS5)[N2FdV(&Ke]UZ_8@DYb-@UDONY>:62a\5P.>cPT;4-gB9T)R[9A=73#]NA]
,\Gb[d?.N0NDUEN;f#Q6Z-VOZ4JaUUT4/FY)7#]c\Rb@Z&&(NTLIAPOT^;Fg)LI&
U<N6Ed32K-<e=/JRKb=bHC16B>bZ(>.c-8^g^1>Q<7@f,HTHHLeY2BZ[>UI\PJ9B
CFY/HF/^HFD^-aW-N[UdfE4VD87X#\Z0_J-9d>\8.M^T,SN]+Tab<K-[<YKB#@gY
=Bf96VBBSM@;Z^#TIVLTC7J2?5B5E4:bI24[[C:06-SVU1YY[c[bc7:=+;Z#Z6/L
7&S,<AW[@?&GW?=LZO9BBLJ+R&7J,=L[V3@+B]bGNM5?)4]e[0bfR5&WEc:7SD6K
49@PZ_U(g:T6_\8?U@[]>D;RO-1\1UFLM:HLCNB/aN#];Zb:;_E&:c0?T@b_S;>#
?(235_NGHXT+^#d>1)_+U)^7XHT3?YO>9OUf-DaFXdTd7aDT(DYXYY75RG9&JF5\
M6Y>35@&,[&=8@W=R-MeGB6:?[7O,=CK#M9eU@TU[;/SNF5&JO-@bf&CPBV\)G:?
9SZ]Q=fG@3I55,,UBC9F9dU,KJYR:C(56>EGKb3J]Aa>LeME)fORV]7ME<X5JZ53
+9G3901X#-?@/X3;OAga<BKSG;5>=.&a(OacS,DL-&bf&bZLS91ZM<a<d5K/6.]R
R&\,H)dSRf<K^Q+e^P5DXBJ9<U;A@5B[&&5Uf\E\+G)\_IDa^-,Ob^CKIe6^IAf]
]D@6gHV/FALCW[HIaKd_fH56:ddU0P]-R/=#f[+EUU)9Y#O25eHe+Fa1)^RJIM?=
KMY5H[\E>6Ad0H70U91LL,-O\D>0FV_UH\DODHeA<_5/.]^RUUW?fbDOF\P6LMM&
[eDSK/G8WY[:91K5QKeZ7Hdf\B+F#MdH]QQfY<We\.bFY1/F;0_b7O2NT&Q21K4P
1d-9(-F5DI<=60Vb59dCH>f&dCb]AE;([ceR[9@J-GH&(b=0V>R)W0ARGZ;ZGTH&
O3/&?:F\bH#IBIEQQN78MOONceC.+AQ;A,6WCA9/N0ZG9gd5URR;E^d-NJ62)=K4
J)M<=SMFYd=_8_^K\+\6gN4YdAYf\(E>XUVJN\QUR-)]+9>LO\90#6#Yg1/gCE<<
1N,O[<E#/fVX9:V0K7?LQTQVJJfT5-Ge4gNRYJ1^bdG63A00WQ5N_H+Y8JC,.d2I
;@2G+,G6:O[P._+8#9B6)N;g<bG3c.<PG-JRW#F8T^)(8K,/LEC9Z@ZX=]A2fX^#
X+BA4Y,S<aDe>GBOK-YbHVCYW@U(OAf)dI<R4PQg#>?OO8.L4adfZYTE+P:3ATJX
cJda+-H=gDbX=O+H]?M1<66YEL.d^3<KL.R>>5:BU#>cA4Z5IM9,E>MYLQC)NfK:
\a.P#\LHAfP+3QBYC_A_9(I2,NJL^;&_@R6@OYReg^AcGFb(&Ec2,R_;J>EXX;Y3
P+X09AI3.JeJT3>U1L@_6HcW<:eaG+X^XGM,O[Z#b,[RXFG,6Q2FDQ95Q#P--1?A
GJC:0HY4@)6VW9?:))FeLIMC8ZB.G\811>&G&=2O)BN=[U.9-ZYKA9,/AU1[Q8CF
5eY+E=N:RDd0&IE,3-,H]A7(L(T,cK_KdfcP7SDf8W=QFWKETPbA/Y(Wd][^)PE8
(QNf(ENI>YJ\ffa;1#c;T3IXO-c<cXZV_G_/L,3@U_4PKI#(=UGaCB9Y6:[W+b6/
K.=cCWgAb?3?-K>3:VcN?Xbe3Q&#;>&A=2W-O\Kf\?:S=#R&X+IJOS[Pd&QD)Y&4
fe0c#1@Od-,M+YVb9A^4?Y9^e4-=^A]GK#Ia\:B(V3G)LV2?:fg@8B9g]ZIZ(YZf
GQ/YTS^3(P,/TUNSg?O>IPH+:<VI)CbUO<IB,.X-Q5e^Zf(K5D8-.T:CM-R>DRQd
.,@+.L@f7/>Q.S8TMFOQ9)7gN#KM=3AOBD@[H;B+3]bU8?U077d4gJT5gSP[E^JZ
#>0?IAAL@#ISfRG:DLX?-2PKG7=X=aSF(H+3a28R-JJ>deS05B@AV=((_>^2J>f+
XD&-/aJ#X>[:XQfNN(8[GP1SNV:ACQ^AcU_@1:bNWA04CSN].>-)Q55b.5<.N][;
@;H[W18SLe#GK>1OD]ag=/8.H^G2UcNO.(=X&41\bJT2O):-Y;9MU4UDUI)<41-L
..;NRgGJ.<OM>BUO?P_5)A=[gX[G.9?M\M+V_A\NY)-4;1F8--9eKggb<D-&:&bT
39V2JR+FP@X#VS[,(6+\W>K,d-_39[67U_a,JaIXJ0Z;a0SSPPOEZ4.S)2MA)K,(
:M:J2&9,EZFT;MX^>((\/d?[BbSd)/f)_eQJI-</Z(>b>>=Ge:NNPBU#_c<]fQGe
8+A(YS]D#;]H99@F)(&XC/U+gaKY5\[MS)d]8cP_DW\d7cJEGABK-gd9[V6EPW8J
gS8\gN7K\DP_DD@0d1KG;d\[H<##RGgCTSLJ5(&(1H()QXfJKLd]3NW,P7CP/_[C
79:6S[b7c,?a(D9Ba)P3E;:Q8PKPfff4dG#6eR<SRL9U^#(C^-C5HFIR6@RA1O_N
:X5L->O82T(g)<1F;ed&21RP,5ea+WCA)[gUP6MMA)WH#AK1M;SZTT:,CH<.RXV&
\e.#2Mf&fe_>)H^08FW/,&/1I?HP6J^[N3:&(WVJ#:@3SY-Sg?6ZB_?YaGg[fY&O
REFC:[<,41Sa:Z>3[d5\(CBR:6+>ZD4NCf?dF830BY<IQ>[/_ZX/bUY:M7TS[dBZ
WF3+&QR3<,H(Q(WEF1IALRXF4O)T^0Xg37LJX/5]UM93SGAfN5gcM9A.C/#Q6ZC/
1X=e@(-Ye>RT<<6Nca)ID8I],9ZD<&[8]PeJQf7b#UMfK^A:;10>b,D^^R..LfTU
D5A0]1V;LVVN(<RgHBV=&SfB7REG@5cbVgcVM7\GGfTJ;6Q&V4LGCZLF[#M;I9#4
0<ABQPJDg4:4eRZ#XHW]IQN6d<].QN=_f+CG3d/T4Z]d/X2].#0d.HbgB#\D>BV-
f0aGT,5f=DWRLfJAAA28)DX^>SI#3Y6KBZ37.IS1d3BBLJU\A/J]<CZPJHffS@<P
8Z8fP[N=:S9B=3fA5TVXKccH88OLfE0>3e5baG<_,VI^9+//]K7CTD1@RcU/&)OE
(P^KQG_6F(=)]MPcEe)+bYRe6]=0b4S>D_3:4bQLSIBM+U+435T4-[<0S;A5>Kbc
]+30;-U+g.7A+(Q1C[;31eIWWLC,TDfH^4A7P[X;8+CBb&+aMAdF@K(P7M;U?YAf
_Mg.HF[a+4Z,&Nc/TX.&2f0JD2\+20;ad7D]9O.,AM;6d(@g[H#.V4)U:^H+b./W
>Nb&aCf.OeWKWfb^-_YZ72cAN:)LA;,NYGGV_E._Me87]MC<+DWU5\T@D+6#6#8D
?Y3=CL\#W1,^)/K1F-I^cN(43GfRS>\F3-XCYS8X,dC,FJE##F;eF[^&_HfH/+fW
Y-Z4J61WG=b]Y4D&KO2=0P)H:@2=8(^?J[9.F8#G?dY6XQ0^F;f@\c<H-=]K)4N8
^0?\XDdcZ;#FNFe2eP).->X[BJ7bRdZ,8d/eBc@9f2RNREg.\9@5#\>)8OH&/(9S
gG4/[C-&B&BU-?5gB59gMbJENHd=3CWE3/57&HFcG.W0#^MH,(f4@M)I>>WEU_,O
M7fTP&VDVFgea[f.6DdU0?,YZ5_#V_79/WDS7>PO7a7ScRXYGRdFDb+;9_J8Q2TD
&0Kdf4)?0(58FH2T\OJGON=S77D2E3E0<C(bD#dSBBeT9KFH?OWbM6^#fHU;8&NO
81SFgM527N?2MFXa\L@aacK.J@^EIXY&)B0U4:9Q,;E^?]\AW^-\+..+Z\=bf;7P
?@P[H3d&YVQ.>Lfd;E;8H=@&CM5DZWXN.=,&fWdc:V],LdWPB^_AYS3.8#CbD(7)
)RWZA(Z/W)@CLbdQg5+-M>-YR@PQE0Wd-MBeRO@+VM8WfPcKU\[])fEDd-<7YLg/
T>M;#VZHcD9-K3CFYX<0(XPZbN@G5Z[J[V]EJV3B-4:]HUge,JOYaMIdZA4g3bf[
==;(XM;A4A95WU^V,#_DWTO@HWL=^8855WO&RXK&?XQAH<AD6\H/A\M7RZBWA,Zd
AFG3T3DdcdE=RZa-V@2/fDKUQLE;A,^CS8CQL1^0gSeaC;)I==d>;1#7e]UEgL&B
YC>d_?#?]8HPLRP[\2B-V#]04XQ<O\QEV)L]dOfIX/O^_aI;G8c\HP5S/,WIM2?]
DWJcRUe&SbP+YI87I#?BTZ_V,QO>SHG^YgT(R1Ud+.GOfXW_,^FA:K+]_@05IPVL
H2/CS7(][\_=HI9?GGQ@MgMfM)F@g?(fU+/5\@-_HZ7\XZ#fD.g1EI6&]&fBg5]<
]9.)TN[7^UMcgC)Q3)[1DWB98?dX:)9cQMfT/SGCP(Kaf5F=2N+#FD.b4.&/AWbQ
:3cV)dS#Y3Lb/b^YK>EcR:6+W9NWZ;N^+/&</12L9,L)?O6b1GAEI4T4I.K)V(6H
KN-a.I?7E]S)c--gIbDX@8J<#9P&>:a>1?\5W0cHGfB51,3]M[>(+:-^BSgTW=4F
M@_UGJ+/42IZ/LP[>PX_A:CFeEGG5N;ae_.+)\D&d8]JLg,_ZKSK\b[@VEYS+=+I
#.B[EgXe,M5RKVAKS9f8@AZbV7[Za]D8A>[/C0>V:<ZUf4?JM&>,gEQ@eBJ;f?AZ
ILT9Iec&\B?<Eg<6(M@YBP\I(]<P1K])(@1)\(4903/H+-0;5dLO9IR,=3D^3=]^
^L=bYWP)BWe?>Y#-/3)eP0:?C,I596P4Ng+7^>3<4/<QCVQJ2ZAO;#(11O=bc-FM
6U/7I_bSg@89X=/[U9MK6S(_.8):?.4b8OVS:;YD[DYb8<Te6Bc32d>XI<F#MA)#
;SJY;SG6L8O[@0f^GbDg?QF<CB^+KeQXY23e4f.d)].A2Z?#PMT65e3R@1P5MKK8
c,8Z4Oa_@&FD[gI<EG?J,URdI9A3OgB?9.(P(TH_6/0616[d77@ac?ZVY,Le&,US
32Y__)#32dc;=]_3f??C+Q:f7259@R0a>Z4S9F7R^&]cEbbOd#K\A?BdYT2E5Q)@
@abNB(_)PZ-)a/BH6I:F@d8eO3FU2D2PFCF_>:#=9:>?VGMO/ZB;&E+@\&Z6[cdP
RR1@(?6O/D)(5FT)5RI=F)0UfX;5(UA#GYX#dX681NQIRd(aS)e-Q8PJY?Og<.8C
RVGVfC]17>c;Y9.0+bO5cTCA@>ZRUG,;:aR@G0HFZ8^Y7;X:#aE@d]d&,&Z1B3C<
T=+BO=@W(+UV?=.]WK5_>cD+8DEY&9PS9);d,5A8;]e;C<W8_JZ&AF>XEKXOB+.[
.?>BJ@529/_7RDfHDdQg/9-5Y2KAcXg\3[b(\3\;;?<K_=\6;801GKY6.,N,D^TC
X;\=P4#=C?N270:\8Lef2D3YB:-\5_;4CLI.-[d/<>4GF^W;N[4,?:)GV&cD=IAb
:4&D;4Bb;^P@8_L;=3-E_/W@[H=KS:YT>]#,SagSU&R6&5C&@6I8P6MOXg/>U>KU
W7G^[VFQ\W30[,H6)C,fd-P83b984@\,DI_0=e(d/@4LCI\]#eF7R?9GTGM5RM7S
(.E3L+0O5<?H681b+1/=E/PEQH?0XD1d?R-5\1)<+f?,@0XMU]\=8+6>8JHX+W62
\8d</V:[aSFGfYA1W->b4)H+2\TNW3;VfbV]N#TFcGd0HHK[::?bWc4eg4H#5^W>
/a7V1]IEbccWC;8S9@ZRc+:2IN<b&WNd6=Q7bN_>bW)@3[NSXLD=.0_b3C9I65^+
EdTQd-Y^afF>RaE]c\N]DF/CZQA8fAPSH07gOKdfQbF^-[:91X?ZL0F75;YB;@N)
8J4L)5(cL7]gRg.+BHHg,60c_dfTSW[IQ/WFebP^/Uff3]#->+O6P(Xc;TU-ZD37
Uf.S>@02Y]6G]ga1&6g=g;#+PUKd8B-/CP1<9Z1Y&6^YWSV#Cf+.>b<;#R)^FTKT
9_dCTY1(M2g38<Y?eH[[<f[#A+RWKY;GL,/cH]P8-1@>\YQ<VI5<.K9c;2BE9<DT
TH@OAUF409Y:_/@_N/a7NUTJ<K13aLN#Qf,E.)d?bg-8DdV78ZVMZ02.dV02dBUD
^<J0MO)cfg4<3_PIE2gaG.=8]HagKSMS3MHY?VKVg9c?9AT\Gd9dPWE<M7=STRef
,PC@aY5d]a25?8+[G6^FbMI&@[GS6gQ+DWE/;/G@V-Q)5JGYf_aXS&O\^@f#+M=Q
PG9,FbX95#4]N]29?D:,C5]QO&-DEZ\WSUWJe=&&cYOVK5K48?=.MTO]AZT1P4D]
F2O8UVC]1gF[+&&I)bQg=,6?(4GaFD\#1#g+2A9<I5ZN\U9H^2^#b,,+DYN:TSXF
^WA8D9K7[[XL;UGBX1HC_I#:?3JeQfCOB,^8X(7?9NVaEO3Hf_N5DTOAGb]U_\U&
4A]4g^c<5[W]V^Aefa[?OM/27E?\QW28[5T(X=;<UE=bUMLEgHH2.a\L+aD2Eb^K
b7;@NNd2F]Wfgg>fK.4;&97BM01^?N-d:L/g>YNI?B_[G]fUW?JJ+,eg@eZfFU#3
CSGO,@=BO<Vg2g8U3#,:;fAc(^7^WTW_0#;Sa<A40DX:Z?WDC&YZGB];\TU7cRHK
J9:WLR)HH^<^?PH)/Z8ZUU;[@WN;0L)ZQ]Z+@bS@795XQb;a-g88<0YVaXMTMZD5
AT&IZ4H[I?-a)=V4GKS0B&M3G]^/0K9=UM4YcC,d4NZ4,d<ef85>,^bgc-F&C8c5
dAA1AD:.;PaUTKN9D7Q#:SS]fL453B,]+Dde^C1TeJE1c<4Od0M8G94EMHLL[LM+
5R<de]_d5cZc#a(cZN)06W@+4:MJGDdgc+QSG6J:@4ZNC..;FVXF4&67/\Q#>;@F
?01f&DOWIaVY()Jeb@Q[8a7XTF_Z6\I9JS3^)NNU4,Ae,L?F66C[=318=?LI<42R
2D/\2#HTVaO4-IRg.@C,WI_K2fg3VI-C/IXaSN^)QPV)N2O>32Z>CP[/,AVNc(1<
XP<H2W;&c:e\VK.9\+cGIgGId6\.@c\?b@)FTU.)^fVGaHLI7YIb<VALL(-GN-:O
[=FQ8]g_NObd[U>fR\:MO?XGJ82eC5_PXSCd#K4b1FKTX71fFC8AEGac/O9Ug^7/
f.bOC<.^-/d0GgN&g9U[aU1a?G)TPK:&74QFBR1@_#A89GP<D(9(]2Y2:;\,dWQ^
@RY:>468b7.f[YLCH)J8V[dBK=<H4D+e>I46QRS]OISLaBEIa+W5.-P-[b1@@=C0
?<FNNU=E<=_.Q<L?=2dSHeQ6T3R,>W8caK<CYNT^Sd?=MT=WgWTG=XRc#E]_?H,=
F5X&ZUY7?MN?0)CZf=\4BL#;&+DCFH#W:YIg&?B\KAP8&/U@gQ,D2NP(6CK,gUHL
(E,8]\?)5AXT[JO-AEb3GUbMT>e_HF04_<OP[VdMZA-I\D:_J0<gE(5-V.N\;g81
(LRXf;\2@AY+<2Q4UJAX.W0G1-;@/OZV\N(;_#@]-fVO6OOea#Ugd2_8VA<19f3+
)f+Mf)\e:a)g.H4\2Z[a?H(Cc,If+f\3C;=^?=CDY)@N7Gd0?J^a+,:X:8PLUW<[
@[8F<67fUfC:E/ee<f=fU=E.3ZXI.6MGU,=e@dTMY]\g669>1Y(.c.7GJR9^f9ND
4gPILT;;7Yd>XRV[-(M])BK9I#Z+cNV@&;A7J\82B<C6_T@107B?1NC>CW;g+#[.
<_F+ZcT;S=dDVdPN+dJJgKPX95/SRgd#2FKN@-U\TcIK/AUH@RJGS_-gQQS.P0D2
6B)g\.^@(5R_[F0J\Z/-S9P7c?T[e4D7:IT0T_JQT9LG075Nd,D:b3\fDM7=/3G:
XK,?/__f0[\,=aV=KY(eXe0,;Y]cO9a<O,E/ObVgHX@8XMNQ;3(S4Fg+?.@U_I(6
F)ZFW;\\<V?g-CW_::Z1_XZJW1Y6:-(/P9:/b4FB^fGcaCgHE0UXA,268C?ONU^F
(/PE]0==R4FS^/T<I?bJ-Z;a(TB/5[SXPLa;?;;WE<>@JZN#GV=eF,P]R(R&T<U\
a[)UR/RYB);NGaeG(Y[8H6K=20^,4#\EN4&cGWVU3b\CT+V@c-^]Q<VgabK>>W>6
CJ<0HeM6IHN>D&OL]XOg3)bR#=La)DW(??a_=O<HD;]45(7a\g>+<2B5P;ZF0b<X
+aRZMI/U+@(aXX?1;8/TI4PYcVJgE&II7((UFL5;B(&W#HKc38F35H9<V[2=N&/g
SHdOeR>20dK70([YMX4F4Oa4TXQUJD&GFdSTb/9U@77#GO=5WS)HL#ZGccK](_UU
K0SV0EA5E9E3GLc>E4J<V-KXGY0HSAC0PCa4F_JWB(_S5FUK]\;B6=Z5J78\G&+R
T>AT;c>10Y,?c.;M\._4eG_7Lf-O(bB#9_[OL,M&\-NBFBRW]9.R4bgQgcd4aR3H
bgc--cR]c.7:gUF4V4</YNU/,ZF9S+_+5YdJPc5(K6Y)b=\J&7gNVCPC9g)aXGM-
VA_Ob\ECNEAV3A1B160BKZ1:VJX0_bFIX2^(^&+cGX+1425B:L.8&.b[-PSPeRI=
-JHb-1:J7CB0S-\\921=3ad#V1U3LE3,;OHR-bF3e&Y04@Q^V#97J4>^B;#Q>0dO
8d6bB:+1)L?\</ET3C:3S:2e6]AgPNMF[@;2d)>0aGQTE,HB\1(0[B&C5RgT]^[[
cM;SYU(c.ZV1B<-&=_VK+PBH&B/A)d8B&&N?Z4:6,19f4;IE5Z^cO+@SS8P:X[UM
#F1;202KS6)&e,+SV?VO&9.8c.0dc;>Af^[V\A_W;fP3_BgLQ>56N0Pf2SEUSF/6
I-D=ff6a0BY<cbcI3<#02:UN;P95BP-c/8/GVJW+Q.X.#V/59##&W2I??bL=7G\.
Q2EbF7>=2BBeJYZ<,J]0+1dCZ.^#]&.b+fgcbef-XVTXHJ6W=&8NJ_fODTW6:OaY
UbI^IJG,A=_RMK+,B/X4<Q<;X04H845?Le#PH^##^6NJNK@eW2GXMG:F@7/W7dXH
O]/+X>)Jd_.Zg:O__9AF.W9VN3<RPgfM)]:Xb,c>S6HQF:YZeDO9W/W[faUMLHU#
Rf1_fMVYf+gZX6<ME1fPfPU_a)e384P89\8Re((QOBfg5:7T??FE],CccF=H^-;+
XS@4OBc#cOOFM1D_KCN)U8QQNN9=J--2IMd(JFNf8#0T;DccJMS^?PDTRCB6=(EG
JbXbPTT:;DLSb6=63:1bR^;1^Z0^G-=I_<<V<ae+(&5U,,d/0M<^P<3J4fRWegLX
Z\^,@,dbc:8]ga.LSSUc</@>C(7?E#U@W<QN,fP9-aNPD:@0:P)e:A-0LN4cYe(<
N9-Q6BeJDZbF_0Mg<69(4Y#f-@@6LB40-2a1#f=_ETU+]UfM?[0B\VeWC64=;Nba
S4=d8\FE:O40]a1T70R61<_1[DGB85WfZB^edK:8T#K99c>Ag7O9gCd;79H3/HH4
Y(FA_f7),(<XW2E//)F]3?&PQbYI,g[@Q5U_@gSWB@+..2cfG<XI6I4H[IUB\ZHD
KK:gW4/aKOE0f7d8:NJd+Q7-SXO+Z7>&EB)<C_8U;1,CKZdAdIR:\K@)ZWCfYS,4
65M=Xd/L<cf8?#V9XGb.&ZU;;=00IdTbM]Xce5?FKHGXEXOR6C@[6;FbAHYF&3g,
dMT[d>=^/-KJ3cdF@G_>F>(D8H2C-JY_RM&,eQB0#a?<CeCFDG]U?I+HHKF/V1/2
Zb-]NbCQ-aDCcSXP2BIA=HQ=V@fA,af]D^YOM,M<#Q-BJ0<<2,ZTUTd5;(PY>1Y6
8H0(HHcg^#&AGW9G.BW<94<55Sg]N8G<0BL27FJGSSHISc?,.VR?OKTJf-8\7eK#
_8B.=EY93R(O];Y_LOcI<c^+2_-T1Y/29NL,RA7NC;#W2bSc09[/A<;L<gJEWY[V
7G+a]]Q7LVTb.Be&E259@WDe@^#1/56WCRe#Na1&eAbe3#+MIWU^U+P)N&]Rb?4U
4e:V)YZ6Hd_EbL[DL-FKaO#dG-PW^F+76[GG<5(O+)adaO>AQ>H7HTeFf9dIURN_
WI?BW<PF;TN6^FFf8gbb[8\05HLad^H&F?R+MX>f>Y&QA.6-OEG]445)cL?^_6Jb
^g7)3;0)[?Y73,GGb>4RKG.a1.UXX-MDGS?g]^I]74B.HP>NIK/5T);R2;#=S3?/
?SB(WHH<cS.U]bDKB_Aa&H@@:FaH(?GJ3=<D(TeGZ4V,H&CfKLQ_<b-<;4W,2bQd
?ZYF80PPOT\QI#U,V@@GAR.M76^=Z4;-Jed))QX?#[O4Q@QHMP/g#F-c[:1G#,dF
1#SEE24G>EA0)[\J+L=?M2+MUHH,NBW-ecMXXaRebLf_O<U]04,?AG@_Va2e=#\b
/-9&#4O;+EYB(/:G[A0HB&P_24&7c[/cCdW-M/1\a]BE/GKSOR7agKD;SVDB90\/
dNE.DASJAEX=WWEM08=L77VSL8G0Af.[6;/DSNT=f3<,D7[4CUR[BTJ;&W1A/P#W
Y.;[&fe=C5NDPc48#=I?Z^XL2<+I=\f_VVW.@EH:Z&&,R08/Y6?N?Hce<>f8A3Hc
926G8TI@EQ7RM=6SL?^FBRHX;.d=_U]N->XRJVSNCd#VEB)Ief5V464B\TC>VR&:
X[@T&_^O(35E-YObCe6+BVS>AV<Q/YI_,eH3a<[G:9656)&#e)6X+\=7A=&+EN#f
&1aTZ93Z0DUb)2D)J(\7769W(eO9@#LELYJ6Bgg5c?cCUgQgXIQ5]g[B05Y[P3IX
-f3QVN-JFdU_\6GKQB\e?ECQ>STAV#W:NWJ#&f)YPBLQ+3B.=Q3U9BZH0D35=K3^
.,;B)QXM]@@KIIJ?(2SA@G:1YNaOXX+Kf[FO_ESCC<5Z0U]f>\f:U[gQU6E0Q)6L
XWQ@[=Q\M[,c]a+1dH#WgJcL.]/BKIGc[;V6U4&]JZbWE&gC0=MFHT\a<-/;/RgS
De&BQJ,M?T]Q+_OfS&(],G4<?d+5OX>T3L^PdgAa]O8YY.aE5PVQV#6Y431U)41.
+BdOYZ@K45eOPNHQUR[+W0MQ0SGG^VdW/<<H^WOIK=4Y)TWd\f)4aB6Y#bM[[g1>
<NHb(<H/G,HMY@9YUUOagO31<?LK^ADE6df:MOL0aWG16/JC?H-K]BA)TU/AV7L>
O[X^)>3cN=(=Z:X-&3Pe<^Mb:U&7MBe(LC,d_DO8)?KHWNL&G:C7\<.7,^+5bQ48
:e[K-/X(-QU3@3+67M&:#ND2E2b^7MS0U&(P,I#]a^Rd,5&YHVKINVe4BERHZ7cU
0c&1G<Z^b[C,MEf^3LG9NU.(27;&,/d2@Z_c8F#&>0aZ<=^P9:CNW+@B3FN26Y&U
;[W.a>5GR9W+IXNIWATEI#H<1bY[UcgOE/_SW>21&>#:FD:L1B4E^]+]I6^#6?DD
N3>+E3[A_8/Y6LT);H4-b8<[Q@d/-3A>V02b[C3LL\A.M-I-7^,X>=cF[1SH](eA
SAK#Lfe&MX_)GK@-;76/X19?Eg,VP?eT)>;fMHBaX.aOT,=(RFK[#,LY=)IQZRZ@
IL[=Wc=c&:=)XM\/7NZL&:UM,7,T+SHR8V+5a(+0],eY_E)/cBVC[[09>]V<Ag@B
A[6:gC\]HXGRcWYVS_9H/749[,>8>]1=O^DS-97.BW;3ADFb#RXOfR5/cI9VFRVa
G3VdF3\A-?X02G\JG2C5]70VGVP2-.f0?2O3TQ=_;JGZ/E557c95\SR\If\Z6dT8
R\:\=H6_=,c>Re<A:,g:7=+04d_<JIT2ffcI]9ZPD9@D1_:^I-9b_WOKD^ZC.TW/
K0/S@U-@RR3&TG62P-+C8I@MSTW]_(+6UBVdZ6?FOSM5?3;BNU&FcW4+78-[GM4I
_CWTZW]P0#+:XL/@Y;D)NFHK@/3[9L<Ka9PbRc?IEV,d>Qd+5/DW:c>7MF,PZOT5
F2@-PeAQEU#]R:H<fL)G8[c<IKIGf/N8AN/<e/7Q25X4UR#+PM0I^g2LY_(QIL5<
0RQ2H]PZbQI^\(L8?VW9De)=OHGc65fGBg9K67g=J4=K.[2I#<bTNL-@F]UO3;O=
&;,??ZHEP7c,9LX.-@f,,;0R?P#3c<]Ra.,W:0_A44]b@,Hc2[OB):#ZGW=?0#Ng
ZMfXV:0Z9HF5?eSQ&=E2+&^)=K/V:MZO+Db]OHC-9YI5I=+LOg(BU998CD;Q7Z(g
56UU^C0CGERPJd).Z?(eIVgdYK2@2b<9HNA]eB&HXQ4N?;2HEM9ZC&;QDeIWP17M
-7Q.0;a4G\e]WJ,2>,NN6;_LJS@<K9>MfKadOA,6=BV6-E/3&9/LTF@=&TI95dB#
B1^C8GaP_+/]&_OR3RR-+NB>^8UgGPcH3I-&5dLFC,/5E(Y.F<AHG-39e-XL7??7
0QZE(IRO?Q9_,A6:e=4g=.QQ3SB?]bWHU;=@/N?8b8H@DF[[K\;fFHe#[M>,.I]6
41#?#S-cO=)c2G46K-J^?-2I6Q;3B3GUG3)O;_V>CI]ICQ8fG5Z&&?fZ&A2MfPHC
(cH.9T6>PIEUM9BQIGAd&V(:9/<f?9OG-e#Q/=31f-&;dW^BB@2f-D.#(PULF>+:
)MDPg_KWcHRIU\&H?1&U6_0TXG.BZ-5Z]S9,OUdY;0)R751KG\4)aZ:9+5JV[3+(
/9^B3P:\0O(AXC=Of@C+3@5?F:JQ@?(<gK=JFZ,8G#GYUY@bf-[KXb\ICLe,F[IB
GKNYJ49UXCD&TW\e6@PfPf2@gZLgc1W7Z>(6gb/TNI)GLNF+2c99(6&-=ZBMGS/Y
3N<cLC.aMLBU5dS5gW6cZHQ>GBLRc7QPfM4Gd[ZgCM^3;X]_V.e/RY;((4D=L<e<
YdN&7#HMCK36DagQ4^VB,Qa/-PI&)?VdL53+I;f>08e+@JGALU(+EB;.T]_(;eX)
=e6eW9M8KDY?bRd,aa+J++]BN-cE[OVLYN?_;/(OF&ZVP8XS]@V2W3/K5K@@JgZ0
HG8cC>^d&0CdRP9]^a(A8WF_8fGSFSGA]c+9U+Hb_WI,fOb38VU(N5Vd]D>Y/CT3
_@(E[)dC:/P#CaTMgA:TV;=#I>.50?@U3@:1I(&&16UXU7HE8:0J:89^/2O^N1(K
JK4WNY03/YJOe6>756G&gKE;9aR)EIBe/RPOS4UD<4,.a>3cegaGM.C4E@UK2;56
6<OZKBFA4)V,(DbHV+C950Ia?K3/GS\Pb=;faCMMc\_a-CDD[4dA;fXg\,?3f:+]
\Od>M+cUA<\<b7)\2)40>ZQ_EI69:6OM2<O/PZeWdK5a\)f8VW+b.8:;@HEb5#eA
d(+>Q65M5?3.B8V4@QJM0Cf8cPPbf=.&-6Kd^&.5?TUfCELD7S_bb\-:=WM0W>F.
;CJ=FeC]0aD_b\Q(6FU(_0gea<+<g,TGe4>&@I8C(FOWd=Y[UT8QKD;>]7]Q41<Q
a,&]<gN)X&dA36V]Y@),G(JG3K]+Wf,9O]<&OMDPY;(-X)aGF#4Z8IO)Pd>7g4d_
E#2)98LdM4M:+5aN)X5TZ3><gIEa8X(L+0U4/;E4;&=D@ST=M(fD+Lb^=11U\,S.
HHN-\_9[285T[BB:.g+VA&Y6,&e\F&0@#QYeE,9@KQ\NKL8#FZY15NgC[L4LccF_
&3=>RD5e2+:ag\fO:0+U5)Mc_\DYRH,\C#cP58HTb//GK\b2Sd9F[=FW[O_C1ZMF
+>L/?04gOOC&SUU^=WDG97d6KESCGF/f=FHXE=B,FRWd>IRB7>f#H_V1C,Fg16?G
L@c=_\\UJ4G_<M-A>5TUMF_R<P5Xec^QTB]VK5Bg]@2LKYG3BRTAZZ8[7#aBdg6I
0I)&AR[+S8IY&)YF)ddHKUHJD9cg;6I0aJ4<I6W)NXe+T0<#>:R6.ER:d3A2Ld7O
Va6N17I^,0<7gNG>:I-495S._+>g&b;914\b0<C8dDJ^G-D&\JGM<K2&A1/]3U]g
5NRGR2Z1=<=TK.Le,CNW?>fY?IPSg@ZR4LC9()/a>0CTMFGDe?RUJ0I2@&[NWca,
G+g5Tg&-Z^R<caK/X[.L-&/1:\QMgUVT@0g7/==RLT-JNR6AL0X=\^P,L:R4dJV6
_bb][dI(8R/c)66_EG2_-H#OdV@\6AO:8W4TE19#G&Y9gT=f[d4#(a68WXEdP\Tg
UWSQU/<)?H4EIb(1QMM,L@g1C)X>b-.&K0-d7HRC656PNS33X^Jb&VR9GHSE>+M#
-]/)7E_;=AfW6cZ6(S33L:_cGFM4Pa2OB?g3C>DBKM3M#9cbN.ZA/[5^:M5[]]eQ
22<D</NJWKDTYf/ZcEVd9Ze\?Qa^+A]NOJ+_Y,:)_Md5RaIfaSNNagVg0_?+LOST
E^cDW+\?1J_OTOf451AcW8_Y2P/R_O?T:+8F/,cg89a,Xa1I/SS[D?]WRTA9P<#g
K0M84&8e^FNR,RSLCcD-cgCgS^W]@A4bGU>0JOE^TfY[KJSafF\7I:EGCcJ>cAPB
??<dLB4^60C8.S\=ec#(KCD=W7;C&)Q+(;I]1.8B=-&eT3^0:LVb+Q_I)D3>HF\Q
XMJSfbOgF)VG2?/.^-7\)6bG<[/d6SFS5(80NgT9OZgXDR0>I-2YNDfUUI/_6>&M
LVUY7Xc#>Z_\]N),T3,XXSg?FBJBG#\2EGOc\</OO3[7S28>GOAFT&4FdFKXbRg-
&NdO+&@YQM</B]#fW.1Y:dF=A;W5GNM4bY7LEYE<_WUaO,fLMAIOM)5O+,=\;//b
H[:7bP>(V2SI8\5/W7)KJ[K_/[RJb<J#T>RJOeU^4c:B+IL0g;/>9-5(>.;N6-/5
?X]L^@?[A#J-2QQe5OSDbN;_-S)f)8R,+E&;(5VY8,0[B[3K9d8.3-:8/=_]^F1<
&>]J]<&&\(PC9P->W2.9Y3@OJCIf6I6aFI.2658GMG/eI@840eY#[3c_G=MMV]O9
Z-)7]OD]5H_00b1#0Z?Gb8#O3V<P8K;;U<U370P031_M-1/D,N,E&@B+@VX?Y@#+
6Hd?).VE]P4_^-N-@Af9,#bY9&fCdHJM+e6/FG5Q?ELNga43g;U6<bCSYZec8?N<
07B2Z.GMC=JaA7bf=-9Sd8N94P7@W3(^GE0afcR77Q5\;51KS(A,<@X[,G&eOX^e
;D[b@,[SK(5=>E+bR&,_F1gLS@d9\QLZ,+Y24Gd0I/+H<R,V3;\I9[XP:>0@e>eH
L2<ZEE?[+2B\)<.dWB=c40\WAP)VPF_PN@f-/+;LHIfHY<]C:PS1bER6@,AMW5X9
ZIg&X]RH4:3K^ed(II6EJUACDK9XQT2OOJYd+Mc_eNbOT-#HIQb53(I?gIR\5b?^
fQWB.-TC-HV)3EQ[b2.#KF^[AS4/J9?/G72);/+9OEI14aaSARJZ+J<-bQ/2-K0R
O1I1&eVD+?8MbNFQZ.cFE4Ld]P?9M9IIeATY=34b7U=>V3M=gOf6E#D3V7B3PMU3
1YgDSd/I;HFHNWcWNUN?YDL4MH<4?H(;,)HBe3Z7@)@J^3YgPb.C8ZcfeQRQMD@/
JSAC3=)>:7Y\ENEVS;^WbK6#CGN3#;KJS649&).[bQYWQTSg]RO4X@;?[/8VPfaS
ZK^1,:E>^E9=08808;L.NDce4A9<4R8/LEMLDH0D\U@_6IUVY0HS0FUbc1TA8])O
d.S^1SI0L,:_/SW@,@[8];3J6(9<36X94:#1YJgW12dGRKL>QG]aQcXSY0QH/H)>
-7/[6J._J)#@fELMEg.3DIcgW::I#&@M-gQ8T3<.]g4),4-5Y<V8?^Y[63#7J(J^
<MS7-Y+=e-K55<EV5L[cI]8()_<9OW&9GLTS;gM.7>FB7-&fXNGfaJFeT_4;NA2=
RZF_J-5\>.G0S[Z8YHAaJc5IXT+5);B\&GN]@BWQ-1FR7Sef=)gbcX75#6e<257Q
9cE8)QJ5<YS,=cPb87gJXJ:c9?]802T@CYL0W7>AJ4=f&;L6X4Og([Mc&C?6\PN]
FUb@LR4]7\+.;^JXfT[,GA]1#H6RWdM?K>X):#MBcbK9-ILHT7XQ_E83)U?HM)<+
:6Z\ID@aYf_.b_]>?0K\4UW^4bE3XQRUIJUHeaLQ\BR#4)T(QQN>&EDQTKV0MHQc
N@^Y8[eeO@VIfRFIFA2-X]^Y-b+/BZ^7E7f2]4>=_gL(_b)A:2#JNXP#;/5a+6_-
2;11/a?NWTe4ZbdU<WC(XVZNgPQJ5UGWX#[W&W&g6f^gNY@0Dg9)R[FDa.F]+@Je
WbBW[e[JfT6Td6IOK[(?^:8C.J>9VcP6/;)684He@b(XE\P.aGJK?_<SD:<.Jd9<
]8.\V2IYYCfMQ;_WW.e+GSEA6//80RLJ((G?\f-[&HP36S4<dE3BMK84e]1e3V]<
8_Ya/U[I:PgQK7W1DY.e(EeW7Ce\g7O.c^X1^NccV5PLdc8^CK9b-9GWYZdBWGb>
^\fJBP>@ADS[/9UB5WX=_\;/+de<W4IVP3TIJ.[,959IL\DcPCB4Saeb]HKGDIF+
&D47L?U(HZ:G9X+BZ0cBaagLgKRb^D8Ue4=J_>.JZ8)1F,6[b>L5L:G&JQJeVLTY
?2:8X05a#(gR[f&T2G?&>gDMRg6ce(Y(C;e@XO)bH[P3>&Y313/TD1//?;RJ5I#O
f-5I@DV4<3QN.KfMM?Z?C3c>DUTJ0DUc?7]5V;&+]2F[75S<U_P]9@+PXU2\@BEa
<_R9L+>dN77L>aU#)M47:ZX?dfGOW,a65+a.;Ya4T@B1D4HIJ[9FZVW?)X++\Ae]
8/]cI=aE^I][U[HG;db-5TZ0F.PESa2W,e5K9C@c1KPA?R<\gX(@O.-Cf^XG)].1
2-PWO+ZX&Hf<SMAGf[?e)OLK/9P_ggf:d8K)]I#ATW_e?P3X+Xc[Cf_X.f9,WOHX
-/b6DcGXI9AM]GVTCW6a:9L^>,f51,U/<abN.4AIe8U8//4A,=ZM1KPN@bg;5YJX
4W=SeV9/Z+KA2>bJE<I<ETAA8Z704M:IE<bFFI0WGLP//..G;eSYe7(=gT3bc5Rb
T_U^.]K.Y?R.S^\^Z>IFg2E:V\Q8,@U[J)Sd]gOB9,FP<DRgVHVVE3(=J$
`endprotected
endmodule


