`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 1000
`define LAT_MIN 100
`endif

module pseudo_DRAM_inst#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/DRAM_inst.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency, 
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:4*64*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 1, DRAM_W_LAT =1, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8191];   // addr from 00000000 to 000203FF

`protected
VaC(fOM0E;XIBObDc<>?_4XCSG)X:=4OKS845g.P4U?D>;YUcdKK1)EF7aX[38eK
/UGb_(g(H--SbURP12(X/WL@#9=BA-4;:#9Z<HI>)HVA=K_E&:]c[\@(Q.730@GM
a62J36K4fK+b8QJ7UJ.bEPSH^a=30M2GLV[X,8,,:AE4F4ZU:4DPb>.3@Y37Wb&Y
8MQREOBEI/ON<Y02;O=R2HS3AH]c46FZEB>K8,1dfOJEcTORP4FVe>>Ra><AF/21
3aRZ,[fJ0F@.KdQ99EA#9O^MQ_1F&]bP)N^O8DLfWc(P[/R@efA8)A.S[2\&+VO0
3_4TO5I(fbKO81-5,I=b7b<OW>8FR8AbVI\0C^E&2\N\<Ha+LC>e1+?Z4XB-(&SL
e.&TJV/BR^N6b,SWcLWVd]DK.aNS0dLPIS-;IX)X7^0TTBPTG=U#F5N519G;gDHC
).L5^E;MC[J/B>9X/10OW;_+,HH)Z\VSZZ;TRZ,;3DMU0B[0\Q@P,Te^/3+7:(->
>QB12FK8=L9U]KDb2=4fAb?RLURc4#>Q8(M3M^><QLd&&-N6@EQG[XA9g\,f@7V&
TABcOK]:[&HM[5eQUe@TdfSCV6VAAV,OMVFbSMY&D-RbXDH:Ic,G82ZCeT2:+UNP
^PUX+U4W(AOF-Hfe<Sg?gaFG_2dSA_W34=VXK8>4E0d-:>Ic#G#12\7&W6++;ec/
?QcED&#K,cfJ@VQ]I:U>,0;L-H+H-dP#>->Zf9->9+gNL@/T@T?X#=dd&,\c^e,G
Ca:[aKXCS]P@-W[0_L3dGa+:J_78_g-gKXYb4,f-Wb<ION+;;IIUF[dVRPL>:7,.
[dH4\e]cVLcJ:OA=1\2(3FIc3C8T5I&[>.<c@(.4\;YE.R]d1P)DHUW@KN.4/2RS
g:ea[^X3c]T])N=<.IFD6/A]c0_>/46,D9.ZDHSN;ZR=:\.0&5;_D1/(5WTW^.BI
^KLV4/=/b;-6F_)dGDB0^@Ea#75#M>1WFKFV73NCb5J^8Qc@SR,3;GLZ&Y:b9cR?
JZ6YP>29.V[eE.PJ1LC(V3L/2/I&dg:ZgNT9<D-eF)ZD9RIO@S)FW9G12B@/B.+#
5TK=eWeOGXR[=U#O6?9XJ]/<.d1YN^Pg//<&c(91cUYEFD)@RfO(.HWOAFYO2&P#
B7P#](_/:7?]^Z892##UJ+^;.,+H(B>9:I)Ze>[Y?_1C8P_+VMOG<a5BLLQZ:0@7
W>f<7d2F.\.&W/GZI=;B7O[QGV=7WcU5&G]-EL?X^R7::Tb9Q37B(.?OSa;4(g8_
BdS_984,b&&=(V>OMM@[AaT6P]:8X@&_4HAJPD8V]Z(,P?7bB,N\P761H>T^B9Cg
U3H=7e?[(,;1N<\9e?I+e6SJJMI@PH6PXDMcX<6)+a_>K]MBVW?_RN-V(/?KJQ.^
CMa@SfN[5M0C\FHPd[;R#7[fX&FUMTae2IL_1&7A&8R?JFFLN>^<-g64__@[S(cY
;_JG.29D&H.T?RM6?NDUT>5&V1H_S97)&cU>--29<(T+NX98N6H-XT#/J1NAK5;I
DN6XeHaaWFQDOM-5XRY(=:TS7Rd(.RW7=^2F)Y.Xae=cbc[^):@VD=3-M[+.O[S_
F1])XaKZN3DeYa_&4eUa_407NHA5&0CJIHZ]BRd>TY:RXLP2RCaSRb,S73G>@&<D
GLZN9,84caTSW;dGF9?>5^(-2FdX[2fJ<:.:ZM/Q\:;5IEIR>6/)?JRB)1QeUUDf
-bA4TED=-bFW_?E2A_f4:ANe^&GM8GfE[a]=9WCL=GNZ/+Jd7N8TU]UU(gJZ^6,E
_LaVL_gH^HOST7N:^]AN71KBEWcb@C3F7(+Ff&5].AaWd\@RLDA]XNPJC7EQ\J6S
R88]QH:Hb-ZL^X^A8++VcJP#8fg3M=XYGZXHb=Z\_2@]G=)\_ee:_L[&XB4;cM)a
1;MK^J9NHJH<E6&_M(,U8=&U_O&bJC90A-6J&O74N\?J4@#_-+2_D(Q.:a=SK>+&
6f:-5AYF9ONLHfaG&7KDN6<X\@G9<>,=Z93fC+.=:K/]ebLbZ]UTc5#&TLc(g2[[
^J&+Xe:gTC;,JZ&3c&:/]EbM\H#\&/5WOWZd@#^<=EDgb2APNf9Z5+W+YeZM<-GW
fP/<1E^ETK)M1f[QNIe:)H^:.CcF3)0a\QZLMPZ;QTe713:=[X6aL(7R9S7[(8/U
7&_>M#A?-AbC1dbZ6ZI(VbZ;VKQ(M1F#OM2^2)<DG^fMB8A:43(T4-bQK4XL:K,g
c#C6/3FM/_GPNG+BH37\HJKHD6EK#A_U<KPL@Y:V@^MR02+EcXgaL>?XB]-I3da7
FZXL&YH/A4]f,3\GBb],CY5LEG)MZ4eR=dCTF3bI:<P?+Pf>T40P2c^+_TCa\G_2
=<0CJ(?^OWdC/JSK4+DSFQ\\8-eH@[.>(IJ:+/WR,Z6N<]f-<V+9Ida0aF2&>+U&
MQ,Ve_CLW6fc8YS.NWCWGY7O^6/5c&1f3JLA=^?FT[ORG>CdfSTe:gZ@CW,?-P.C
60TMJV\BbR\NNFPgdKP-^PcJPg.PI,W#70X&5>=\9P_e3/J99O^J[TV^QI#8-4G/
]V=PDeIRa344>U/.H)F-=2FYc5Q):7C,6A?b@#bP(8;(HW3JUe^b]cfD\[f_Sb:M
U.XgSRR^TPa;gK;@^g[G<Gf6CT8_@UVEX;fVOA[:.8=;d;0cX#\+HB9d]bB<H1E;
=[NMb[-5M[8HS0K[R?YVA0g0Od\?#X>@+RZb(S(AfDaSW_/b2[:-A>4Y?,X<V5>J
aIDXQ3Z4daLd6>X839AH;U/VWd6FX485G0<RP/1NMV>UQ._K@IYYY.PIT]HB42SA
1OZd3>9/T:-dRX4Gff4^AX?Y+K?95FLf;OGJMO\GG+EdSA(+DD:GZgZR:O/(a4W/
RfU^]Z,g^&fLX^:4GU@d9PgZWW1UHL:O^IcT[O9Z]YTc0b.U5EPBNd?-W7B]4GOI
c^^?B+?]W&\d;HZHJ1bJXG4T_9PSVUDRSI?2U1>ZFS2K)]aMQ\]7K>0J_,351N?d
[@K8I5T_g.(UHP+HCH;d81?XAc_Ac+c;_fEISN06@#c8&I>Q<_H)#C@6-\e31G]/
a7fO_.VE(eZS#T0J(9(I(D/a;&/[\DT,K+[3HeB4[I(V#/@Ubc\9Ed/^eHB;Q_G4
gYA;V]EI:CccJ._bg<.DAA=66K-^/[6VJ.^+X7N&J;\V&(<XKC&.:gF48>K>UPJ3
&aM/#[&;HN+g;9.Q.9P0LEg)HEY@LeaeC.TA_J10)G@WbM<?4KZ@G^/RP+B+W0,3
\5(Wf#de?N2[+fV/0]NE[ALNG@=:#AAK6+K;aZ9YIFAcF,?-<[-(AO\;OY?-)U<+
/Z<Tg2A=AP@JDHCN/aV<db9EbDV.3YO(K)&OG:@)84IAHMf7@b\C@U<W.39GSA=g
6a&f>9;9TeG\/Se?3+fcf\)LEAE[\\#)],eTBQC,E0@F7#T<@/@D<a,9^&Z5dZDS
TWDe8XWN+/R12(D0G<XPWN/?Ob#b1SJ._aH9fDHa4>PX>L8(7eQT5LT=P2K^((E2
N?=Lb38L7Qfd00U2@@M(4>MJE?;9b20Q/3ELb6F?1<YX0&FT^Z::Q&fX/URIR1XF
Of6OA_J8SNNa+4]DI+SAd0,LC,&8=IGMDM.GHA.ITB=9//Y6cVGJ_V<FOaJ(bcQf
4FQgEPfGf-U9XNQ9d49?/4P)RSWCX/Y;f,I/)M+^gF5X8fT)0LPOV^I=V7CXaU-V
>;A>A=:>2GQ?.0>D,b]bM7V)17A>>O1D][eG98]LA4\<\:0<a[b0(ZHRC&\_<\D1
_3V+P7T8H@M^R=HJO[)Q_^Lff[#GJF9B(2K/R=c8:V;Q@9_J#fYH;0D652UG,aHC
Tg6<,GG?0MT5IbT57LZ9e(3>WWQUfcT_MULTC>ebA?_P+a=S<PO4+ZUY&AO81UNN
6P-X?4e=+30\CeOJ41c=S>-ID<8=55^Df.N(_-;Z^cD@&/\d5,X\XUegYWGgO-JK
adbecX^3F>eN<MZH,fM<);F3;dJ5M/##efUX3\aQ20PX9UFP6(@6RTEcG;=/dTR#
P#&N>]N-\-;[Tcb<MDP>;B7cN]=APTTO74W43W_D6\ECc8B4.7c1GB)aH];BA(D4
d&DdJ6fLAAdWF/CV:OK7S=P:A.BV,[3,(H:55J0>JK\_gAPJXRN.a1A2]\5V.N;K
F0da@T[eO]<\@;V@^,,&I8cR^O/?[KMEQ&GMO9L<e]Qa&==D\7:5J&M-<be5bHLE
IgZ)KSO)I-QdeIJb]C#U;>&#I,PP.DV-^6-19U-4:X&.e9cL;>\F-#>SSRa/<7BA
#P_+fK6V]>(^+bZG<R[QY4d^JER79-#A\Q8NA7Y<d1d,?4Q9fe2XP>aL9CERWDX9
[+)0Ge>ELSOGJcW23DX=._7>SDU+]e0Xg3I(Z.(K31NM.XCJJXZJf]1=I0;\KScG
V-eLX:(^G+[b#3D7ZYA]6f4CT3U8N#Y5aE8_FQfBW7g)^IV),=g4?<#dX2C5(^91
4__9V_KaMV081&JJJZ,M#;b.3A1Ba_EYYMBR=>Ed0S4G-EGfWN2[+MIM;6BNL<YO
4L9:#>5JW\b7QfPgIV@DgO\.a#(B09eSggR>S<BbFb.H4>b1GbXfd6)3L[aAg<Ig
]@L5HM4-e92_9QI24WH/V=RD<,;(<ROYeU?B.<-L]MJd8W6;Y_7ESO<8dCWXTEQA
=NbJF2J?HXdXZ\06A_g8E8JZEc0\YP_cA+&d?A(&18d\EX@@JHZ&8^,JRI+B6C5,
@g].SfeTCB&J:egaa.3_:_ET_A#b.PTAa3<BT(.]G+MI[>;32FH[2-gaP?BKcCIB
5Z9K\R<^fC/Z0a-OX--?06IT7FXV2dQeUQ=N,_I=#dH;KSW<[>-0d]D:98#B+R?0
+6ZUHP;5)Z@P[;Rg5a->a?bbWU.FCAG7YT&71@aT0X0-NFS\:+9)4-ADFJ1=I4L7
U5<0Wd3S_J3RWD>PXT4dA@b&[&#\0A),K)60JfF++abaN&?5fA/BAUIOKZ+CM/1O
Y;\DTRBD9dK-S);Hg^<M4P3/[;9)&egaGE33_6:L29O;Cg>B\9fHR7[O_7_E;P?J
0D^=JfK0W_#WH.F2.?_@fL5Ob/3/P\ZI6&JReGK(Q/_.Kd.&QY6JHG<),OSdZ,;&
G@L;XNWT:W)KO3W9&<eI]XfW:G<M.=afGA)_8e9KO-M7=0?Q#/1QI&AD([XZ8O)9
Nb>&V)P:YZWOdX206c[KE2dQW/RW1J,-W[DCI5&8K5.T95GB>Ga-]<[>eIEQ6eKZ
;]OLD4G=E46HV]E5BMQbR[E<b:8Y/g(^gI2BK)MS#;)eeEX?Tb#U[->00VfB3-40
M-eQB-^J5YXA)E@f@,()aZH?6X[R04C,Y>E\Hc+])-f+2H,/W_W\3OAY[<A&_]H,
IN+=H6dQYPZ-P,DF0EQLe1K7_<dGK>@4R3QE5LCN+d:MF6;3dR?(L,4&]YTd[O;1
gJRO4UI+CCg6[ZJ&\AF)0J=;G/cHJ(5N_-F1H\<)#3eF8^F/CdNVbac(R]_9,Vg(
,>W-/=c7IF[eOUTf(>N-/VH+E78W&I_#T_8NVB83=Y?EID#C8L#f9\C3YD^GWGFb
>B?J005YP::;aPbAU<_.,4UO8M?_/YI<\4/[(;U&3]3MS\8UXb5,9OJ7JaWF?.J+
V\O+FT>&^.)CFQ/e3Se)[GMG6G\f@G?I4AeOe:ML^[/L,\IBB4IZ[U9N3(K\M27I
c9RE+?:R+>40_JeDFK[fDR17/#C@A=N]O@ZHe9ff;;d/+gUfAO([</6c[WX?5H:=
WC<2@@V6IS#8R6=c3K>.e_CPUF012:6Xd0#BWA7P)P+1d7e^5N\Z;GGdYF=VN.fQ
W./,cY(YEaC^#U/f(<ccKQ,ZLP1J_D]24eDL[d4P1#aVH?QZ0K\T.FJ,K?eZGc-,
&@dZM=3PPAX-GcB4>cGZ=G8BgEK#=C7ACH.)D;c-NX(^21SLU1QTDgbJPJA)UNN:
^JRgEU0#[6UU2cd<[RGB=fK(Ke_P1VdO9@_g31^,.&K-L&EWV/3EdB889)(4:@II
\?A&dEUMU<60dZ)8(]#?W<gPZM@[,ab>52ZUfDYHAL+Ve:.:?^.<D.]Dd_MGdDVG
;0\e3dd_OP6V4<=4V71cU_N[Y[F/>G;)GV<[S=DG2.aTTNLS3,/J50EQB1)>P..]
?/YT.?IC\+Z/#<c43A717,\XfE:KH&DM3LR+OL1\W9gC[Y1QJZ@Dg3\+d+2Y1f<M
FHd^EA(8[BJKa;bBAf)L196E3/gd&_fe_(XC9d:T5XO+?Bg+>\0&a/_07J,FKYGK
4I^aMV,/Z1O]092<&;(cC;03B3@;.7=<9V#5G#+17W[g5Q8cKZIc[e]:CW>=MWG#
1\VDFRQ-^b0([bT[7,ZTSe0D-0FFV]4:0)+b4+(Zb\171B#Bg,T=aHY@Ycbe\dE1
>PACNFS.&S>KV6[WG/.YM@U9[,(C--,+6g+BDVe2N=-FbI_@NX4N3NFCd0e1/ePe
NGVA)A7D=9:.T^B&cRXV32VKZ^P;I-AVfXMR7Cb&;89XF[g.O/#Y(TC:(d-a,OC.
?d)>4_SL:M-7E)I=<BUe7a7g9^TQW5MBU-EU)YR-Z)_@OYb1K<[R+.\)Kd#:b=U/
4WKf1X@91/LHZ,I(@L51Q][8/DPPK]:ZBI,@SV3,GYaF=V(#9YEg1A(W_cKG05&-
3c8WfZ((S=00Y)9.\,THC11bQC^P[K2>SZc?>_(WK1MFLKY@__Y8U2aUC:GU,(5-
:S_#>?I9_+R8d5_>409Z5=1>EPc8?NTOCF->NcHY6YE\_=d>,7F>TNN(2MSaY)(X
S._+eg3R1^T/WQgf:+O@b(4c8D8;T34TZg0+,@MI7@SK=SHE,aGG9-USJ,HWV<)L
dGDb^KJBSXA=/f2@S/I4I;6Y+LAEFU-#K6M9I4Q07+G<W()Z^-W0RC:]5EcYX)2D
1^2?[_=:,M(AL9N#H&-;eg;K=YZP#8<cZ3W554[V,=)+PQV(=c]62Y23+MF>-ebY
I?=UP>W,8/EJfSE_?H9S)D]WKIP344S&59f:Hfg^1Jg7gF1d>N047TA>IY#4S__>
P?M8S0<fgT/4DH3)aJA69aTY9f+W-a,Z;&[>-Q+W#)9(SLL&.KCF(Dc<#(9--H?c
X5;B7,1([B[J<3gY>QL_QG].cf=4.[]J=W_/XDf2J(7:-&09\W1+:QL&X^V[]#WR
Vd8GYg??,@2=TfAQ.PeIdPFL)Z5RBMPag37BO;.I?TD-<UI0IA+>M3O#WeZPSfOL
1\c.ZS73a0T]#gBb64FWWG1OK81[U9,6A@>?aD<^Z=b;+-[B@0f[-3D)WP:KCV._
.Xc.W5]7BZE_RZI1PI.e8Ta.L-CE,C^^:+;TZDP(INBcdE>R00bVdLEZN/5@Yc\]
cKD5;^@>3R]b;=NSOYWV)cL6UY/C+02fb3.IFQZ67_)_D^70a?8b&0g4=^bdT_Y/
D]B\(+&)JU2V-cOW):D[HBa97?,/4=E,Q;-(53@;V#6=QK;-fD7MJUVa:I<<W)GY
F9+1_RTK@b)T_2d:Q]8-EfOUFGM_=Q;JLV#Wdcc)FdbNCPaeXG(359]VcRbA^YEN
H>FK-Q@FKEGK2IE9E++]#LRId<b6^4D,;V;Z&XIbWQUB+H+\D[Z-BW&8VbY6&bD0
I&Y/;/ON=TZJL4@5DU31_6(BWRN(^XbCb;bJgFOa(-I951&,S;)6CT.R^d-cXK>K
<+-d?SXgKRH=2OV-;_FC3WFgEP6^4J\#3LZ/:-]PNa[@+,P,EP#/&XB[dA\0.=G7
5I6A(.SC6TQC(ZUe7-[LP6-G30WH0MB3MIKfAJHYE5ac_>d7T?D3gN3Y/Fa2?>0+
R>N[0VY\,KM]f6TE9-#VOU:=Mg)QaOZI5L6Q@6#.N9^V0P8UIQ,<fLCd3_Tfd1?g
IAf&dR?M7I2cY5]Pb\bYXc=GB6O]0DX;\B<1(0W6[71A648-NTIAGb/XJYL4&CD0
&XE<LR_#IA:gP3(8Q.CdfNU0QHb<,g3dMLE,Sf?WV(_)Y(2W.GcO-_9HbA0:U6)U
F#Z9@-AKFVX+XVTA=]0;/O>1=IT<Y+1W8^80e_aHW,:BQ[J)b;?9^&C@/?+gHXQU
@P8[2:.D]@fGD+\A]5;:A;_:R6U41C4&32@[+F[Q)F7H5YeIE,d)@Jb4M;aUP?5>
LWP4<WN3L#f.K^_d=Ecb<-YL8/B9\eL+5B^CM0e1f>]1CR3[E]=(\-99SK5fe]EF
HWOG<)ccMM&<3fZa78GfKO1OXaeg=NdFC9928[]5#4_AJ=AF;NR8gU7BLFf)]T-C
2fP__^Y3MBC:HUBZ>#QgNAP[V0]4fSZC^P;E[MJCUdR(>,23J#gD?X&a1JeAA=Y6
+-.+5SKL35bVB7@2HAO?:Yc+=ZM2fO>cE^PHII\P?egXUOOg]XbF:Z]4-8;):A1F
A::>XBR]Hd36??GeU]FPYKVb:_0>P-1N?SP(#)RFceS/].@LZ+EG/HIVKJNQ.B+1
P-A64?XV_:?YJV+aaB/+U)O\CY9>V)447D;F>:3DgO;^[c^M^\,M?KgA(gRB3:C/
.D3<dC-VD06V0B158aK9fE=#gDE4(=4/dZ(Ug/7KN/+cA#:b+]6aC55J?@dR0+EG
@C[>U7b4Jd-+CKEg1SU:2CE<(a#<d6?2a>@ePKT&34ON]0NS/R[^N6+GL\aH+[FH
=7ER-]+BP;&B3:Q,:M4eJ-Bae8E3AAJG?KYZIHLN;KTQ,HYD0S.b?e^8]6ZebBfJ
fGaCT7;J_dCFcJZS#XP6U/7/2,@6&d1B(&=;O_X2,K.U#F6I7/:O>8Z?-?]84,)J
bccf8+a,W]ZG8gKAOS:C(GHAKMFegc7A4)OX7dIMHXD/b23U&e?dMW\d#BIbMRb8
]7+a)]dfUX)COeO2b]@4cE?788ZZXZ,=6TeFg#JHa1^A4VEI:;HS&,(VBT6->NfS
7Y]<&/H[gO<;J&;cg7_HVAFJ>#0WD6:,)R;Da:g639TGU1Sd0&?0BI&&1>LIBH:B
faDPF8Be4AgK]>7@N-WC&2^6c(a??Z(V_bReg.-TN?)9GOR08UA54<WL]_5.BTfZ
IK_+E0AZ/JJ>B?\&#<:\WX/e[gK5-#XFUgH-32O.;7:IaKH2B>84)&,S&JMV5#UL
5&/<JWIBJP+YNQT+2TLCg0JU,8N^b_-=_^d8Pb0KCWA-\[>N<]@RKd@J?SO1]6]Z
(cX.#aQV=CZbg-A#\E^e4BR<Q#b_1Ub&TYbgQ(CB;B?/UHUK2,WC-4ZNDQXFcK8V
Q4TH44-ICZU[&.c_1B8fP]7(3cPMV7Td?O;FWX#PDGK2K:=__/7)>;0aZ8BUPUAb
246XHe/#a2@\A[6S<I6KNQ+9gPOc/JT2DK,O-&>1G(M>a1a<263#R8(L9H;-/O74
a[N6Z\S4.Zb=T1EW@R7:-ED1)(HR0bb&b5#^(Y\&6.)d>X,fF5\2fVODXIeS/QOY
.+9OISNe45<GfSgFSA0A?L;([U+1N09J1M#W>N.bEF66cgC/:_b.Z:#/fA@+WQ9U
+^7fb2_2]HCY27XT#WeLW7cV)B(bC)NP^TS0XF@ZD^DDMTFAIO;cGBAC=(Q6M]G^
NEQf0#=a7<)F\BUPJHRa(7Sa\d^E5YKI^c.SW9:\G@)=8X??GdKVc)W,G)T5W/dM
3Q[HCP??NI>M.5bD7D(I8E?gG?USB1FO9>f,Bb_RDJAF@PE7?374F4794:4#Qb>#
HBT?H<JQ4#YO>OZ=&af#8HS]g(C0;AF@bHA7-JAKE^:]]38BZQ>^]dWa1Qe1_W:b
a8G->/@<a9c#FGRCB2^0I[(>;8>6>GGTQ(RJ+=^&RY(2J9@K?bc\Aad;agg;H[JW
[]^PSHVD]Mc0>3<_))2GU?gCe&GS<:+IKIWe]GT2PC;2UQ]@6E(\-THg\cfO[c-E
8K/@WBN:c^&LKe+FD4e_c5#?)^8^9eNTbDT&49(g[5BS?26c8MQ04\D2GC/TO-N8
S2.@5-;)F#bTCB.fe-YP<c(DC3U;NM7U##ADWZ1)PKHbfFaIAK[F@UQ<<KTVIOUa
c>AC)Q,b/YJ___=E2G9YCNKYPDgY:.+76>LZ&aT#Ya8QG+\bV;R3B#PYK2K9c509
FI+Yb2PR6Y7^T.WCQ5RFbg9E>9V94(M(NTYK&;EAa^=_4bW2Dc968U_N0KUN,Xe#
KJ^K<1##85DbK-5V17DD-F_0Z?N9Kg&YaZ=fW/;WT7U:UCIf(]>_9=R/?IYGNdB4
P@PH:?L?DL[Hfd.(ZI#9Y,?8EDX@B?Z)e@G6Lg4M0;TE@^beL<KX#XS>>UIfZ7<H
(a:VM2-:a?@C-QD+g]0\NF+;g>)5]V+5DAM-fKDQ6@f6D9&J5KcQ:71LK9W7>GPf
GJ03@ZAS@a?fAH,)N?XcUZ6/&ES((.9AdY=OFfU<&0L_Y(fB[VOYOWHcGF3fC)(R
Cb0Hf@MNL6FDDa[FeF1,K6bM<T[0H1[RQ/K<]ZG?eI0Z6ROYPMfNWKJMM,U0@=>=
8+KF>e49Dd-;,SaPKK/7,E2AS2@gGVY4MW7=2)^97:;IG5\ZKe^L/>)MgN=1DBIQ
HQ(>JU8>71@[2BEJ63UOEfcW4&>28],ED+Ed4;=9RNbZ>ZM=I/c:117XUQI;#-HW
-VX^=eO&g/Q.7bc/O4((]42K<WeZ;_,4\:g,37-M5URZ6Z#UgT]6P8E8C20QPd2W
_;ZP??(cPLJB4c?SB3U]^FXE2(0#PW+#[#AEG8E-Wf;^ERFQVLUS#,NV]F97D6&G
(\5#-U#8^H(_[>V7LU,,\U>,J6/e-W7^=C7;^SL.ZWN4;O/IgC:,5^HgHC8/2.++
N&(3/6KH9QM@Z^Q^aJgf=3HT=P2b1JM9-\#cMVPJVg._MA)R7FTDUT8BfZcN5R0,
QRRO4GSM891K4<;bIg?D&^Q:O,M<_(gLPQ;N+=:S_)e9Z^<N7X=]?Q_6Ee_,=VSP
YIX.<A)aUg>b5X8]L^]6Rg)WSN<3.OJU<H,JSc37BSb,@AAOU0O8YZ\:5=BTf72A
?^))]D,bE?dL[M<#EO?M\CQec[2+.<ce2Fa5CLS;c_^1T:>YM:SR4YF8&b>eIN&S
VF2C[#7Y2#fQ_2LZge6FCcfUC=0_Z/7N4B\88_AI,71)LA;94cT&JeUAS0\&KOQ:
;/.3-\F@4S_^B:\?g^H?b;@_2EZ>918NG9_g,.[]46:X+B5HcLF?81/&W?HaeY25
Q-&d@N2&;_eUV,#8bL,P>A&#<KV4Q;0FC,Z>.&85WS[e]#50-5=^DCd,@N&2UTYN
[>(I(7-?-PdWdf_Z>JCfHN06JG99,T.?C53PB+F#[+<]d-G]@L-4,^M_=g6c+=[+
C9?faLJHWA&bIF(CUK-aDB>0:=I9__c#QebbJcQTR7V9&eDaZFbd7CHZAK)_5UdX
VB.^C5?TV3/XKEE9++Zf-_-JS6\X6:&W;6]0fJ_c+TW?.NA&,QSKSd7]VagGU,Cg
eQg3ATe@/K7E^P_LKATcddI_M96^\6^#=(<Q.AZ#89U4V3(]4e8ZKOdUQeV<?A?X
DHW>+0W@gY(&2DG<fA:W;6TRPRKQReHc;5P+>A:K@ZE?HD:4<.BC:O_8E@Ff4#X]
4)T&I#a/\R4b0QO0:XW].fE/Gf]?<821gUIbXM<dPLMWS&Z8=[b)f&0:[LZZ51_&
Rf^SMN<[P0dVPKD@=(bQH#8/BLZdOHW]dI,@6P_b3P-aY..3Ma^1=cLG3;U8PM_8
7g0ZJ[HcLU?;/E\?W?BJQ^dE#];X[6X_(I<Vf41?H=>7V77;&6RJY/J(E2R@4&fK
bL[94@,U5c/ZTU&d21,\?_5d^H)#PYPca0:V16(a4^,1.B?#E9]=;Kb7M[IbNY_6
d2UX?DVD7_.Lcc4;VbD/PNb)3-_PDUU#JFCYF6HNLfHfX3VCRQS2?&dSHU^C9c4b
fHYdb_?<g:]gd^aEVZ;O==2K^[&N@PM0S05FLWOP?8HD6EGbPWT)J:?8(0gd.U;.
:(TFf[;f3/g[8#XD][XB>ZfL#);5H?eTZ)1c[V6HI]89J<f.@ARfS(c1<\3:#6dN
8)^7C@:K7I4E)X&Y&6O@eIS@cK-W[ML3?XA773A4;60b+>F^B;UB)]M24Y\#)FRg
9VT\P>JQgW>TAd\+YI?DN&2OI80-R)[&7gEB33JW1K=3P>YR_b<;b7]KTI=>A&00
e6PQe-_2:Y6O_JM:@RIY?dV9eUbS,VgC2I5<Igc]dO73(d3:38IP^5:\+@=/BeKa
I2AEPM315eJ0IQ>7&ZNg&@GCa-_7_/<ZGdMQb/;6<\)\A;68.9:<&2U8_<_[IdIU
<GM#[ISA@CE&F-=GJZWG-^HCY+,V5@@IKDW<+KGdN@]A06L9HBTQ8@[)+99VSAPS
R[;)E7QB[DPC0I\^a/S0U6A+2EE68aK2gJ>D/7Q&=BDF0E=M]A6@(C#f9+LgQSB7
8.7>a7g+SE7;.RaEZ\?P5dEFQ7#Q#>9V4;J]Bd3Q.(_M?R2NTb8C&QcO111OaP;:
C/HPRU)Z5LccER347KX4ba)YD=D?WVF?JV0Z7[5&.HYfPS-Z,5@@GRfGK[1B^Qe5
eLIMVB8EcVFNIF(WFB)]])N-=IX]F]cTLJcL-EdN0cW2(9IQTcEQX<0?FWN-O#:5
=TF\N3gMZe/\f8#&[RE)#?@8c64#NT?B_6/,1@Hc;_NW4?[^+8.b#G3SI>2P:4e8
/+(2OXec]6-OEHT-:3TYa(J2T[a)Q>VVKAZacUPXM9MUQ+FI&N&?^ID,bOY4HT=J
M8R\S^(JZ=(KC59Y6eTL/4]fJ:RU.E.\]Ja:@Z\Rb72Z]Q9O<RP+N21E&=eOIMb\
PcLMg36KXXA=E;M#/d0d-^3)-ZM9bS1G)6b+=d./bI-E.#JK.?7]]P]cDTE)E>4Y
71=:.B(9G2eLIJ-b9+fMJ_f(W5AV]TP\)fE\&=;c5[,P3ddJ58L9,N-bI[JXK4,b
gd?F6J6W-KP820_8>3.;+=._7NQLd@)4a7b7bS::S1=<+/UPMb/4J<H/MIO78N5R
f:GJ).#;[;&e:HfcT;/a/SV9V40+a;+K0@9]OB5b1(ARVEYDc[5YPLNOe]]WDa5a
(XcX>3/KSI3ZBOJbK-VVF@))>R(JRQM[U;77-2W)X(QOB9]K;B.2Y_\4+/XcC&4K
&TR]=(_CCWc97ScQZXW935UM[7bd]H9,[2EGQXMg0(\6(380A&:DbZgWf7=T64H\
b_9cb[.IP;N1\bI>PJf+PKTf4(I1.MK;A8^#M-:A\Tb3P(;\e1R&gB8?UJI_d?5A
3#e_-MX/HB&LI]C0g@4:P.SIV]4Fa\LJO_W^\d<U)CU#W&J5TS8SCEF3;&+YW>X7
Qaa8;>-=43GTW5[_c@;-+E/:4I61cfS)7N73(8?^=LQ-f_bX:^K6I:O]0-9VB<8O
9:)A-I_;[IZ27C;54fWDL/@JDdZ[eD8aQIWYDE&)E#-&9ETE9,de6RIcY#b8DC(&
G/BNC^UC;FeSE50<ga1EO\f_ZH2:5CKRXG2(Kd(e88J89dXbV/QV=I1BEK^:O@VE
?2&=GbL+-N2MZ2[FX[>PMJaSQ6?1ZDGXCF1H3b_R4#R;Z]cO1ZGLL,3..71c>Wb_
Y8H6\KG<1RVKJ5N2V([4+2;.MKAB6:^?d9_+6&TUMWV-&@J2Q>d++f7V2Ug)M7<+
X?ZZS9RE_><>R=QG<)D3@FZ:=g,/)-K<20OC?,/c#agD,c;]f6O.E05e,MI[1,aJ
Nf3<_X[JFKf@6R,cdJ?@Y/]-ANS(Y(gGcLMfOS5S,gO9[SS>PK3<X::ELZP->[4:
fg,&C8]#;UHZ.B/P+?#L)1Lbf.FDfH>bf\:AZX.PDSA1^13a>aD^E@Z446FW5+Wf
LQEb46Ie\^9B[faUP[Y<YggALG.DcI:,N^OAFTAR1?D2Y4Sc&+d^_AcNWBKLES/X
Hd3FL;1b]1.M(Q->ULdX@YN^a^&-V]E&86#W3CY0<CUMB,DG39JCOcc+C.T1L0O0
+)-(R2./Ce8/]ZX0PEOTK)9d2G]F;#1;#YK&]KU5)A;2E5>JgJ5gcKAI),BGQ4Na
gNPH/(+^,.#)\0I=.)E#2[-UC2MZ?4VC<7I1+6c55TGI@/\JF[2(=OF=3,-ZW.cN
:FP#N8Y1/7D)SX++^#Bd<J=QL25&\)<A/4JFgYR,1YDGcO96?+@[L7C(Xf7.2XcE
^VX3&)BK]P-7<fa@ATcf0-^@Ea@_9AdbSMH.+A]4>YSL<Rb.eX8CMa^P3VRHPU<_
8RT2J.D63EdIC9KYGE7T64(YQ5F8WXF0T5&I1-@M:^W6V1J/1^6P]YIMX4#L\egZ
8^)[f6Xc8=EO6C@N\EU.QK(Ud9)fg5E?S(>@-OMf[3-T.J(]),;3H3cQVOCe^8a/
X4H3>M2#W=H14YH8YL/cDgBCdX:(_BZK1A0IGcG@Z3CK<d(6;b(S)M6adP.VCZKC
1I4<Y6H+<VKME8)b31bZ3L;2=Og,BA2NT?>NPUY#Ig.5XX6]=Y_XT05GZ?1]L].#
)g3^=#1.TEU)-I5NFIAb&M>gVL3&->b?R-Y?63P<7E:-P@EPI1YQ?03bB8ZOVEWf
c?GfG)5YacZ6:J36P&3VaX53_NMFbYF]^PBg?88f=8R0JMfJVOR@A-:KbY#7,(>H
,DabT[_+,91-78Q65E^FKe#QeE8:RRK:@?F#QVROYRc1=OK_@,?Qgc6OQY(.@4)e
#.L,<X8Q74[]UE_K<3DCJd9P=>>NP&LBHJXda+0SKXDBbFe4S;J\3.H)Pe2Z0#-C
aPg5\/SPBgQ6O?G1Z(FBc.G_c8,U1CLXQSd3:/\e>ALfPW^]BEXUQ>SU,J2QF9I;
7/5[Rc3HZP[,JV[FJOVeM_(_9^P:cMc].g_J)B/3V-]#+P&L=S^c]aO+ZK_X2-3E
[#YD(.<d_gK0@@5<KYc-WA/&W_cQQ0:d5)B83dS3b\SZL_(ec77g]9ee+g)VIG<A
54=6eO.Vf-(df@3DW7\&_XYJ.aP];6B_U8gQdE02A2NQ4DB3aef<;&_2S[Ae5&D[
S1NfH5ALf<9Tc;c^K_F:Jebc7JcF_;6C71LIBZJWd#7D^AaDb&1;&@I)O2cOVB3M
?M8GcZb)./+Y#+R0N(>D(4LEJ-cM<^CH_:4bW<Y9-gDc0.L<AKHf^#<GL6>,@95Q
dd:YXS/-VT^g#R/^_d_82RYY/.TDX@;a_EKc>9^Dc,)+D-M:d/@eO\MKSWB6G3d]
TeEIbe\fOF^9;65W-]<TT9PHNgESeG>Q3L\T14W=bg(faGNGO=IC64G&b++_Qd&b
gX#?b9:?M[7Wa,5QK?X\3I:Se>#fC0;TXKD-]J&Zga2Q1B9YN2[:0bAA/37[[QEN
Y?bW?=+9PBc1:G=K.beDUc.FM(U]L+NF2^NU;g&Q)5;3YA.a,&gbO;.G<ZbQCBb9
:6&V;8CF_/>2?(]&aMTJ6,2/<WGU[c7LW6MXMJR,d]SM3>P(e/U08_.>//dKg205
H_V=FeFf;5.7/85SW6#X&VTY5;V,H<0NTV/T@gAW(:\VH&1X=_&e;UTfb0\.P1@_
V(,A;_OFG]+\VX8c#I&J33-0B.\/>./B#&PK4J)AO]FJPU?\1A>EU9[8OX<a4J8/
-ZPQ9B#UeDPGNg>PH/-D,<T&Y9+NaGBD^WKO/)TdH:bYJdaHGe2N18#P1QRcaMM6
O_9eCYXXXB.GTeeDJ2T@cII6;P39THR=X8?+EG3f&9FU)W4Q)<+?OFDQ:]YeRW#;
/2CUPYOaRDP#URd[fdKL,aAW/Yg)6U?_3ZQ)KZ4BUY_D,<JFO@GG\aI.22=HabEN
?HW2]UE\5Y<E\c09C\3#0R]628DVB2SS]XTeDeK0I?eM@Ea4NKM@/)cE(R@A_[]J
+LbM^8eMgEf.Y_<Ic]1_0),L,Y19de+?3:dL5DI8L_dL<])5_-57eO@=),X_,E^X
N@;.)-+9>;Q_JEd6I-aY=fC:e)LZB47?=OJ0S-TZ+\cd^1-G(O4gBBc[F3)?QTeL
\8Y6VdDH==&AYBPQXQc>)G>aN^99#HQTZGa-29\8fKSgC&;CA_?4+OXRP/ZX7I6#
:DcP<g11S<9a\d,_R#<3Wd,Kb^L\:3PNF,DT833#]^b1f7/#J#-U5<XQ;.Qg?1NH
;UR=W@J;OSHI:^;f=,&B,:SGQe8:/;J/O(B4+UIJ2Na\0?)+451+4F)MHX:VEQO\
\-WgK?NFQ4LD/g<=729E3XHNK/XN0P/YB4SF:@FgDe4EZEgV0I)OdROaI=YBB-=B
K5SM)_L7[O:O9QLWYG:H.,eS/5\\Z=eJ3bF_5OO/T9Q>,Te,_H#f70M143gT^PFR
38>.cAUVC?IEg...ARY&cMa/#ZC;,-PHZ+(H8c>5DVY]7Z;[A4]0U@g\)FY@12.P
V692>;[R\P#1_U72IYGT\3&V8?,[OBF54]KM7^V(8I3a?EdAO98?.?0O:EU:JZIJ
(WLb:VI=+7TNad#/.@?([3X?1WM/H=+KYQ3J_A-=ZG>5c)[V0=733XL6;18>KbR&
;RPC&AL4/6F-W>=9((Z=aeSA^;@ON^+?OO9_eYbgI[K=585K1HHH?,R\GT&]=\>9
eK9KF2\Rf(A[Ee272.T&cZ4.VRP9S@7Wd.e1<-.)GYQ8&FcN.I^NEKdR,Q<E<Xec
YHfZ6HKa.C\B\\5<D,V26EU&IV9eBf7b@UWGQV26HdN(R+0:O8B4(VY(0Fa10+&H
8F]YW&VZF5U[I2-:CAL,?G_R7c9D)-c0>MdF=?LOV\>BSgPE-/Q0)@\14-:_(G,5
()&YXcJ5Q@ObSb09^6c_^^=1fKcH6-)#O[LQPHOK[?(#eTMQ12<@B8,7K.=(F(MQ
(gZ^NG>OY,7F=Z&=,_LGON+-ceUN4G]d1O1+8N4bT\1QgA.A>^.cQNTd@]G+T-O>
c[,c(,63cF[#-=YTG4=ME(6V&TW=IA&6Q;30F)cQ]:Z8C\@0)D(dI<HIQ3A\Y]_e
47&=N1-97Z-X]]GTQ8Za9J-1ePaUU;;_M(@6=Q&g0[c0/VZ/d]8Rdf@RfN\FL/c_
]SS,]aK]a7+#P23Q=He/S,EB.HGES2feGMQQ+aAcN:6D)?DO5-5FQKS67-(KbQ:&
)f.S\bT\<+T?Hcc-W]G&,Y3b,/A:N)TA]4170#fQdF].Y3^?(.TQS0a8:2-_,b2.
7#[\eXO=X[ASFbBfS_/>]48Y&<bQ/XgQ,6-)&cAK\38QK1,8N]E@aZ];:R03&50H
LJ)J;b:4>K8J)\YMd)J8&\?0W&Yb:T?b-:]Q)DbMCDbTbg+d[+=]F\fT?NGMe9;3
9&D:5G&6/@T.#]W(HAb7f+.6W>V8#].>/LT7F^eXYbHX,NV#O/PS?\,3gYQ4E[\;
2A-a<9e5HX@FDc8d[M@ZRZT^\IX\=RA1X7eP2;]V3X@Td@=6J-;27XNJ>UeTA/+0
(?+8/I895;Z@9LVILRQK_W2&C.U(dIZ:/HRVR]1<^7?e(Kd^F+#K.5/J@C:d24?G
Fd-T]L^a6dI5L@e&=APP0^Y383,967:Hb=@QE13;Yg^AYHL7D<SNY,1\PaR>?G3V
05AC,9HY7e8NC?FA+Q,29=&]0]Y^N=4&1cP[3\E5</C))Q54V.G:.FSZMdF^W=@N
06FRVb]@>^HK(^5M]GC.[>;4^&/GCeR)Z1_S]TNP4+/NaYR4g+A,EONaB^JJFJL8
.?/&.>eS4=YX(<U;V-F;C/LQTX4B)b.5Q1dLK[E/\V/VgE-=?-WOV-e6@JDCM.>9
gg:\gQQ2E_04\MRQ^e_;:6XN?cPcY\(#YRETG]FPF?QY&YK)H\+;5<ggE7DN?^S[
3&8dG9K7FXbBK^-baF278S7)I>L.P^(/CVI6-A41:FELNc[+-L&LaQ3?VD#\)QQ#
/^MI]&ZYf=?gO1A,SGT>J^(F+RVTL#;[IG,f^E+Z?Y(102Z3bU2W#aF]af83;TGG
0aS0?;RA+<<a>O8]J=40E^I?BMZ?Pa9BU=<P[V3c5DHCCBG/:+84.^&=)P/L-GK?
?8CNCNcOOD?JC/&Q^Te_&.:D+-LHg9BaOM=)8>0F>C(4YObF2W;W)f4B;A>A/Y@_
9W<5TM5S6G+Rd=UZU+UZ709=b69/O==4ZPc82P&Z]KF,N/Z\]C9(_X.d19eC+D9V
\H87[0cMcdB8a/We/@G6UF-@;d6>7TUBDITQ8b&dI>[B[&]-7W_1W:3Lc<[T1@]A
8eN[_fXWA<:<T2bcDc0d[95ZF6>KW]>NZIUXMY[g,F8;U,Ac(=\K8_4GXbSXL:^,
9)Sf7-cZQS3O7dY/cX.UbgQN41/G,1+WPb)A>_.20Z0>3O.Fb]2^)2]2)b@5S=OV
OQL<6I_OT[B,<A6GF=TEebJH1#S]RK\_f7OP[Nc15b=?82>B=\V:CT2<3:f?g7]N
faC-T9[F^E);RX3e7dZ:G5_]:,9UHgF?6bcBGEIOWZP3\/U.5C#S:NW9W@?LR<V,
Qa7&O2]=)<fb@0#YXZ;LJHV2G:f#8f=E08FgVd1QA(;0AZ:W[QEQc8)(1MO.ObgK
4ab@D0a7_J92P:Y&gQY]]?LBYR)52BUeNdY\g;?FJNR^UD#<LcLC/>+g_1EVT,:^
K93LET0?B9T_@</fY9KQQ#RN(Ib>d1:?O);M(5;L>_Q-Q[GK9-W_)Y=(0[XX;2O<
7Y6RgK<^E:c?SR2?3UWecGJB/J2GITcO.^<\;07=H9FZ8@&I^/b=e,:Bb_[E017O
3[H&ZMfV#d<a>OGN=1AZ;dH.33+JX2a\BB@O+f#]Hf1P]:ZR2&B7Z:GdJKF>L06N
[76OIC+&GOJfgQL&9LIVg,AeB\T7\WLGP[:)PIJW3)c)=28WI,@?/[-(HD)KQg7J
(O=9-\7<4BBZNQ<8--TZa]JT4b-4@T^#T=#c(&BK(f.9@JaC]EH=[@eZKP?Gaa_E
UZf8[MZ::S95b]E2g/QN>D\0MbWea4JH3@Y>RaVGbFR9J<>fN=BPc)^]].49==Q/
AeA=C3L;AT7b/a[,FY&N,RC>KL=)KF&V?E\M5#b3GF4?ceeM2DeGA^dISJ(:\FaY
1>J;acN,E0^]HL6/._W8e/5I.7Y3d:5MOFSeeM>^d3-U1L9>YH<d#Y:0H=5/+XQV
4/+I,2g^d2\WF.O[/?M=JPK62@]_0/RY+.>6Q5CZ.KZQF65M9<C4>AQ:M#A2ZeBd
3^JVC5PJgaLA?=8-1:HQ_\ISd[39[GBSL?Bd51GDGE:8ATGC<]9f7Og\g[2K[e-=
CdG;+?a#B8H4^V^H_^Ldgb[IHB+RUA/5TY\&+2g1@9f-8J;&BUc)UW0JS0,R(.+1
ZG5BP9HP3OSPVUW?J/JgT7RMFU7.[Cc9C2De^bI)J2c>AQZZYW#I)1,MG0HAK=PD
_Dfag:B2CV_f1&<Y_CDG/acM?2TU8N?C\<[D/C/eZ3+G5B#-5O@CQ)U.0,_MCY8a
aZFWVV@gR6K]HY-)_;5S4=&S7K6?3EM5W\M39<A\B>F8Ec>+/c,(.[d[6?W(=egC
:5P,Pb/97K4f27-XZF7,QDb[e@6fKQ7\^O:CAd+>_:,HE?M0#KGNG.<Z:)8X<g3Z
dT/PCJ?],P]RfSb-e=,D[?5[+;5U+9,T8&<?#A,5aY(S\X&BWU1c93M)SZMMX[93
B_-Nd]6L(.9Jf?T5]..FIJg#YcBP3BAC5WV..#2=\B-9II^CbgQ0CQ>GJ<ETf:^T
Ee#cFT_F_B28CS4-_ONHDgZH3cD.d-CA5cTGAfd5F4GX1ZC(L2@[-WR>PDDPU#;4
K@3JTA3#SBF]F_K#4aI/3dP87WbN?5X2+)L7FYI3aWFg=WL_e]>FE7MGPHPR5+.T
U;#e0\7U\ZC^9Y/&bCEMbJ3XM=;X;H\X349^a[0)M?L9ae=/Y>Z;>4M0D10@4-G+
I:dc\27-HX34O@X#U#&f#\TG>LBK04_I?EZ1@6AE1g+:U)[ag#a66HXF/LSS52PJ
-C5ED51&=91]6\S5\PE1>3fed.UM>&fa.9)P>,F04e.(1C@H>Y4@7dBC>AMH@4=&
:PF7#K7^)V81dFQEJ##gc#cM/:V=O)V)DJB7A^\Ccc4,L]1PQ:8U0T(6?WJ@H8dW
]?W5X\bV6C[<8bUAZS+#6_E]O.V;81/#caP^VI10gYQ1\]P23FUY)7c.>#(LMUX;
@YfODF]PH1CQ-LbH;1-_7F_7UVY.G5#@[)XOR,1Z)6g0)/8g_c6G&FD1-19=>)II
F=YU3I8V9ET@/6;MPdXU4Z5VEO(b(F7XPE_E24SRaZ9NWM&5>WB&JF^I[7@F6#D2
=5e-BJQPG:S.XMZd]T@=,)IB,a?:+[,T5>JU.gD(0TET4G8HDaKQUSV)d\f;19/G
@4BPCVPb4:aNUaJ69AWB+AZge)VP[gE\,a107?0d_<T=G;PI+V:e/H5DJ43[<eP>
IXV?I,=;:/f5)gcb@E#GS3]C7b5&^g6XGPB@6I(a7P=Z<TaLE3SfGDZ1gRUaJLcC
>&?R([EXN<RKZ=379=cSXb(,Q13^0,72L_(bCIMB]VGA4/QNY=IZ#L4?YXRRE4.Q
6Ha=^X^&^6V19R<]13<H+@KA9G9e[GIE#4&?\8V3=BG96U<3>aPM0gLK(#,M];G_
^ZH?=a79C]aP[Kg38<?@afcc1Tc<7_)?_QH&#??b5a-X1O:8b#QD;:d6<T.S&:T^
/fME01Rd#7S-AJHa06;e2Z.3b_+#F+Q=K:D]F&-SA1<J8g5V])\K0]a]g5IL[(+X
O[?VR0Gb(/BV0aS=2_R)2#f7eX>;>4/._a4Y&B6QMA=.J\IdFVaN45D+XA(F=JPA
6C@?W5\[_K@c:W8F5=5=0-?bB#4d<?6A6;D[g>FZJ-X5DGg5Y-^O)gY?BZIA/?Me
-;MWJ.H5NF\gA[g77\8.e1f<E<?7Q1SU,a4aX8F=gCQ&[=fZcdGOI&]HO0be_78E
^J61Y.+N^L_P,8#&F)gc4M7QAEP28QD=7K)]WE0NHX?:T&HJI?8+Md&XPN3YYIcR
e_3H:>@+/+[3<\bD?[>Sb6G5N.44_5bD>D^K3>1R+>(@/@OOZLIP[I_,-c+IAPPg
f#b(PFVHUT=VN4C>?N4671/JHg<+Y=S3Ug,>CH#Egd[<DQe.8V3_U?GGIDbQFFC/
WAgQ1[].].gRU48OH6V-6(A)??(BXNDCS(b.7F;#3<N0XaMTI8bHD/#e0;VXEGFS
2.&=B=LWTCb3;V.PT-6bH86?>Y::9?\DY9VbSbP?;;4+,=W3T6Ig^)4_^1B&,BAZ
3b-U35IN2K_75BHY393_+B<-<2>B121W<g3T>G_IM#10=X+DL?F>D<]K>,:0,41?
BZ96>KGXdL5T1K]Pe8I[6AV4cZ\757+@ZAWNR^1[98bMIAONSX;GL00g(#geD)RP
2/<=MEF4H-S06da/G02+@=\F,)BN(A2R?^X,a>^b5NG1BRW_RPcIJ\-/XH>)R?K[
\8@GWNKK3T^.G2SS?U>_O#RGg),.RXM^C@(>W5D+N7YDf]-:VOQ8aB];ag=])0&F
DV1Y(U.6PP+(FFEfUY6dZ>E=]PL4[@,P88#[1>IZOO)28^O(R;E1BaY40?PD=d=N
9N/12.T90OGAU)fe3A1E^),#[)B+:W=7+5:776JbfY^PDN^M(^RRCYK8K1:UG.;,
W2KZ?^9V;,Rd+^EdB/4I0E51Y4H@<gF+11C627<Q>W>Q/&O11@LJA6;T]/BRRdCa
f1-EC5I9SH?(WVN>&,TE5(c[)DP,CA)/>K[K4>G+LD;03/8+<\8bPGU@IXZE63WX
,T;\&e]c+I:<UHSg97Lbg&G+1WM+EbFbVH?<LZ]QO6<>QUS.6_O5Q?c3<6M/WPI@
Ha#-N2fP#+6JR<T1)_7M,Q?E2D5V/KYH1Pc.SW6FUPQ3eD^8Z>(L8>#XONBYP:<.
&:b,PH,Y:Ic.7:/YBf^ggQK-QYK7g6LLN@aFI)2U@);[OB#@3cIKK-(8_3eg-9L-
FdIRfS0LZX2Sa@J2(HW^9@NcE)4&cbgT.D9;(5,B1Ga1UfEHFYBKe])\C7C7\_37
<H?NeX5AD,LV@145GH_T&X)&T#IX,J?,57g1[50f/eVbddN193FIf#d>\?,NeA>@
^7L6B&8OMCVc;N;+-F]8R)R0M>P+bLcPKL1U#&]QKR4TUeW6URK^+<9cb_T+\fLQ
ON<U<0>F)511^WFTI,>D&MX>\B2cf(WV2Z-W=1;_XMc1H<0>W,CMKQgXGEK]d=P\
\8+UE^?@T2P=ZTeGPVL_Y#?f?3\eRfFYEV@YT6<eIX9QR[,Zc/C:+)f/8661X=X;
J?^@WXZb<c-YINIHR:Y92:LM5c4Q@Je.+g(>?^;EG0)C\#AZV7C=IR>e&S3C]B/F
\ZfRCaAM2[c#2Y_5PHO45+O8_;PCfM+IeB=9RA2)YNUdO5ePS83K.4.=-;d;7[F]
(\(5LeGYQ5TG2_Z;S<&7B\YKKIc4(O<.d)MS@>&<=Hg-3C7(FQSE&Y\^Z1[4H(&X
NHDA/<J(O?6a_;R71_&\TUS]<\F_=IPGNMP5Be-eW)5E[-UL_AX9<DC:O5H#A,#C
5fSFSIeaUCOc5;3;ZI_>\Q#+)VR]A&5gA^O8aMMc-R42g0Ma(;;2OSXKVON/dS:Z
R<O2OZO3bg>+J3J4[XFWA<d&/Y&@>,F]Oc?Zc+e4Z9)@B_Z4f-;))UP#\W=ZKA9c
@/fMJ6P>0+3?dD\;Dcf9WbN])AX\]P[3?a-#bJD<9)NO1X9FXU;175OU5YNGc;I_
1?Eabe_VXZ=N8E;B2ET/N-[,&QHbeCUO&bJP4X=Z9I[Q#JbO]IDgWPdI@05\HaZ4
S-A0M7E725c#TNVJ\aU\Y(8&S[=cQ.[\KGW:\YAAdcQ]JV2)^c+bb,V@.<CI7S)#
J5Z)/2fG8OYEM-Vg?/9^:L<OQV)-)IaC33.SNgC]/6[D8N1H3Q(XgB\UO_#d;U14
ZHHSN9a;S_BTTP[<EV:X8),:[?2(QDf4\K,W3&C^F)]GC74BSIDWW5fN]9@FI2Yg
=,I0Ha/TC6BSLd0R)7:->H+;;>]C;V+/U>USc2BTFdHdV-\,MQ^-g/THO+CK<V<6
?fa[1dJ,5#@P>R]#Q(+f.5CLWMFYS_LV:aXD1g(P34O&/X5-A,McI:gM>(SgHg1O
\&-/_4]b=K#?G1XJ\Mc^C3?gTE37OOT199UJXGCL_2A0KOMa3KAZ0)KF[Z69-V;9
GD#U+D8@C_NbCRLOK3<A;b^O>f./U10ZE0If]ggHM&#a_\&K<K(@[Q:0FB3F7>#L
5B-1EHLI?f;(IJgQ>K&47J9,Oa6cdQGOg#_:-3SR@Gd#O(+F@_?N,_8[YGJYS(3D
T2JD=I6B[N7.JR3_)QOUBK^=3f0eI@;)X>b.0J[d/):PS..=-Cb>c16EU5e(b+eH
+Q.9[cC;\W@;X:>fWST^\NR&<8NG_HL[BI3[5+R]K2-4[f-@P=TQD:RNRI.AINF2
MA4Ic4AI[FG@3cggeIVK\NTQW4B,ZE>1KIAF:TW<1<Oe)X^SX@/NNL=:4_,[WMJ_
#6?V@1AII/J47;W+].GII1\],J5VR1/b+Sb(O@d.a[HeB$
`endprotected
