//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2023 ICLAB Fall Course
//   Lab03      : BRIDGE
//   Author     : Ting-Yu Chang
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : pseudo_SD.v
//   Module Name : pseudo_SD
//   Release version : v1.0 (Release Date: Sep-2023)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module pseudo_SD
`protected
8deHMGL:2dH]/@-8f.=+MbX2(?V)CV85L]\UaP9&da.&)\aB9BA_()+V^,1&[.+Y
/8B@PU^II,#1\;_=9e_c?bA,W,7S8b;C7)5C&bSL[5;(YRQM[cB/41cS0NdeVBbf
453.BNJRKLHPWS:A6XFcMYgJ?\V\FH+4\fD/ZcJ&e0H,U?c?^RRcaZVPTEbT]:)Z
]PgH@(6+(P2@S>>Ga#9IbWFZAABNL(DP1c<G;#+[2-Oc__XfRO<]bFK,eX2M5A>]
B\Rc1ecVbHI@_;V3O7Y7.GLGK47]a3@6R?)UN[Be2E8+f@/0KXG;((4bbW>H;W7N
bI0_KK=cg7_B[(\<#J0#=f0G5Q40O9O)_8=/QM8R,d5O9>d)L;K?f5e/?)ZdgDL>
)_fK3aI.[d1F=CB4S,Q60YADLC+M0Gb_BD#S4[K#91G,EC[0SF3R&Q7#9(]_/fG6
8KRHJ+ZIgO\[GQ0VVW+OYX?91eQQ-4NCE:J9-C]4A?OP#+XfH#[L-+bH886FMD.O
cCL@L.&-=H#D<7]>WD/@aK13)=f>45^eP,\@XNZ>=)0.a.a=&-H;GK+#XTZd4d]c
GV@Kd3>QCOdfLZ1O8]c,Y/g0H93,)fBdGP(#J5K+_bR>SPZ/QE5SG[J26Y039ff?
Pa2[^B#7S:L-J=DI.Z2-Q-/WL)@[G8]eW5Tc.W6)JX^ZT()F[9cN^T(\D&dDQ9P<
>#2PU0_-,E;+?1Ye\;2:4I18VRc7W7SBN\EK2Gaf5V9Q^JIX\T8:JS+Rf[a#L#ad
&U=AKK3RF)S\d0=3T\)R=+::Q&6./7fEbM\WRAg,0CJPH4[#=[YM@Z:I\N+CLW3D
T^,5W-)WEgNePb&M4/[FWc>F2@BPaPU4AV-eVNb)/1&dZ,cO)1RSZKVc[/_T5634
O+b]gc4#HSGR[8P>HQVBUSe:&#WCT=Y.8T_5[[23\6U2XS@8O1e1^(.<f/,9S5>:
310^4MYYffEAGWD3ceO43P204<03>DD(GR.+0]]TX.H7/AM^GcIa.U:W6,6(VcU_
0J0_]59H5(c:\IA2_5aZ9ZK?(EAaC9]HS?IU.7.??F[UZW\Y1UdZc/Y=\[f;+:X9
=].1TU]g4Z)=b)?b>XL+(L+#KL,26DPaVG5?:HcFa9+f8J8Kef##^NCVWL_3/-EJ
#X:JIU-H)-aSZEA,K<W:3I-C::fMGX^#XONg2W+?M,\1(@R50SdQE6SZ]2<HRO#Q
(MELU8/LS6H@]4LeJW,HK2=?U_AfDTf<b;VR>7edA,LCUTd3Xb2<;96A6BFA3WJH
SPB#HC0G4)fR#<-=DDWfSeQDF<>F2e#\JQ_C3MT4-c^\(K>D#HO^g;^gD.?UZEAN
(^K04J^]cGG5SUBT4JI0I[3=2EJQNWN#1O@a/:N>JNcRd,;0DUFK.cR-<6/RA(V^
&1EbW.:R#,80gRKIG8Q1:LZATe:@E^2#@6:#J:J@K.Xf_M4)&HL4(ObIKS/>H:N-
_LWC56KfH=c_<d/?S4S\GV6Q=UI1BOG9)[g0FU_E0>CR&/JeJ)[1BO4>&H#V\GHG
[,Q&FKZ3?83Q&I;;2+)-XFZ/&b4-V>Zb?ARg667+,Ue<4@[\YZZ8c/gYLPI?E>:R
9=#D.NPY&P#_:d+AQKMeWB8[cF<g7/#Z>f4+>7V)WO776-E8=)KMW#D^NZW8P<OH
HL:G++=KKS/OHJ.8Y+.3MEfd3P\Sg8JZ@0WRY>e4BX_ZD;A@W3#1FEfWRQV^5HO6
1C/A@K=7ZgB;6S#FaSd8I+0E-Q15<OA[6dE;aV4(L?MZJG3]f]-RNZD:\F@dJ(Od
g2_>C/:N4/LJ+Jd]39:P][2AG,>D3<^;d?CYPI>X#II;?6YaQN8LH>XB^]4E^>,6
4J7&7+=_>I[BFKH).^)1UN?.EW&J(:+010QM3d\+>IG?MHIOI,f/2RTEb/\M1A4]
\5,/dM+-DH8XfH9:CcK[#5IQ2&2),W[B9CV(=5aW,,8cc\B;4N3Wc=aNXH(OMaZY
ccWGaL)L.g6G@T-=5;g<K&=g(eJ#K&gJQf8OBL7TR/d^+6gGJQ7b=f9)(OTU34Ee
AAS+5?(U2X9)XM8QZ9KVe>Q?&,FfU;\W<NA?F9g^7c9dR[@V,46)=#-7(g0[cD5B
AA_J_B?0S)fE#+EKM-/@QZI=LHe71bF6DL_URgW0I;W+-Wa3(_P]+,WaP1J<2WFO
Q/:/WCgc2D0#Y,b]1eNH-4SA/6LDE1Cg,9@@GX?T=b/<<AAa(01F=K6[:4I1D>CK
UZ84V)(0:fF&.D)5_eN1K#bCOGYbWL=d)I.N^)OW[&R)U&7Z:BQ\Y&Q::X1-_([5
IXCCaQ(.8@Ma=1[E\5<f\PeH8T(?LT#,M191g46Q4g@QN)Y[WY+e/bW/<ED]45<g
FD6_+V9E]BK+=YCEgdZ][3^C0RK#A_&31g4H9H9^;ZU4<:d7AJd],3#<_S(S)>g&
9be)5LA^Lc]S_Ae.R\R6Y/KO1,<EB4F-A)4c&^,(c9KKRB&ST=19Ia,-Fb\<U/?\
Ca:#Lf;PP[<)?+BA\QAXaVK70XHAW[OVM8?41A+bFNAZUW7H-DA]KNR3fD=6ZHdP
_X\.Gg/_DcG2,9GbSDS8Y4S2OK\XQWS](5POPC+#M/MDF-^Wa8b,bM9:B\IeZ/AZ
=#1_4YYL(]DXe&Z[8Ef\,TaHVcJ:FD<B)_B-WZ;@Q2IRNEYN44M.XHASN2N2bTIZ
R7&gBO_Za:\c2\D,58Q@GXI2Ga=XA<fF?5]L<H,^Wc6E.PG3[UeF,Z?3d?<(U]Q-
26cO?@:IZE8>QY8KY<X</8OQ49_gE.;S_)>d[bI1c&-48B@N\D-57.K5G87^XMVX
^O2)NW;\4;F<dF)JK]e]P2SgF0MNW];.VSVBZWBTX-LKg(bde[+<(8Y@TJ/8_KBN
cT)F)Vgf(a]aVGgREeQ)W<,A,:6-IW9NZG?/:PC5D4+RcP)a85S;T^WF1GB/:JVY
6M\b.)a[M#2<OAS(:c\_OVO)4Kc3)fU9RL[Uf3;b5Y.^=g]6>IZIE@X,d/UAP20F
G^HeF>@_-[]RWVF3JBT>9+X9]dFA>GMO(I5.>^BFF0.NNe4[V##015SAc^ZGS]S;
V[H65/DaYW8N3@+,.Cd7.GF1UJPAS:KP^02W0.B4DKX+_cAL-P(e0X?GBP;L2QWI
85^Nfa?+XgYeBH2BD2)=U\GNJ3;WVR^b<bJgQ=&b[(.C/FNDa.)b:5<R-JK7Y]_-
)FU-5JS?A0S9W&N<b+Kc/:_HY@4R1FG#WU1<9&?\)3/d_M?bU>M5E;K>KFN\\:gc
=HK6(>deg1,D<KMYQ\C1HZI.TGEDG/=CcP6((13^<,;,ad;//bg^05VTP1JX=CB_
d?C,:G88MRfH8eG/XBD-7TC&1E.<d,ZA^eDcECf?B04U134G9<ILY_#];_b90+>>
N@;g>&D623#\Q=@L],B]V&4(Jd435H=_4[3,^O==169=9DD<6\U/14OXEUJ=9gFX
GRCNUV8@E&ELB(b4[+[K+D)VccaM0?(;.\U+Z1()-&Z_\V,gCVNB2(EHM?&6Fd()
T[?:1>=-Q.E7:P>:T+Y<IW_[=1df4ZC82EUIb@W?Y3=Pb)b(RK8OWDF?T];YM1A]
V5K]>5Rg-#?A4c^cD)db-D45CLS>6MbCbGI<EJ8R^PcI@2a-NX@6R[=VMF/O,TUc
;(4(WXd.;\cIZ9[c]aKTf)E^gW4CAgI(KLL39QbNPaJQ#+BLS:F)1e]CA<>M]^aK
\L+VD6[.b?D>>K\RUC[Fa[dd=,d0aI23cS7]32S-[45(:cb;,)[)-S.Q9M9>XE<)
,c.4E:4QMTa8aB#_]56M&-+F&W^A#<KePQ>#4BIT/QNS6[/KdN;^d[W:E3&-G_/&
.]81Z-#8fFQ6,eUD1g/a2FKZ)8FBC3a@O-+d?#A@[a3ZDdHI;#d^]e<\_AHU:0LN
BKD3S11Q4(&g6G&X(_3<Y26[bSeS4;<.^]O[]OWHGP&CN,EeaQg:++8;K5N(LK5B
Qg5SYGA)3X)/-B2/C9U1V@a6d>SE&NSP+]+deRA)R/#e&gQ31e(C]#N6XZ->@,5^
[DE#8bD/?O;LK3_aG8(KN=:e0&=K0X9.AEB_X=+HRa#cD9.UI,6a-AJ&b4RN=CAH
?Y-C2MS;);;,Fd??>HTA=E]A)ZO2dWLgX=NOZ2K:AMC3[&XWfF&(Eg2;d1aaWU1\
=aQ^8bNNTLMYf;gf[:SC()bC-O5\,^=N3AWLQ9V+,;-#X(<#WUXY9G1_^)YT,FC;
PJ@]9+;=Ag+7L/=ffaI:g+Ic+_EI_A^QdSD,CPK]1VM8@PGL[EBeA[]0B;?<T0WV
;Z,3Z(O8(BMPB=/.SdY09S)3Z>[D)b[I@0Z@]Pd8B8B8)O:E_gWY(),68d/KaB7[
dR:ZF:2N]OP(5QM.I&]O?b+:UEc\Z,V]eACaG]7IM3WWUdP;P9ae3^&EC66Ed?0_
&bYX\1D;NdV^>\40g[2>+0DT?d;B=fH^EZ7cEAURGC>34dd<W?WQK0-\Wb_6IXGA
HVT2cgG(X35VfV_<B/27#NF@RB[@COT7dH^RV0QHHY.\H4B@TRFV9QcYIVJTbTf<
+?>6gZ>@-3<e:5O8;XCFTOb>>(I3/dP-KPcK;eSZ:Y)A_2DG(=_]&ZR&bAE??ROG
P+V^cRbX&)B84Z\g1PC-KgALdbffR[SA\;bggZGXI(K\c<,LA&S+HIU7UTC6M#--
(&RX3-f=,ZJAMIG>URYO+80>]Y^Z]OYN<2B7A4YA-MBHab.@,XPdaa3=DB:8]6Z4
8>+[Y]2TO9(:9XNe&Hf5f^DeIV@W.>@8YIQZ9c\?,CQ]Z)C4<e&+&Zb1Y<:;)MB?
5_Vd+Ud1=+JQJR24/O,#2[f,FO\MeU@)dH=gS]:G.6dC/00;6U8fg.5MC.FO37c5
/MHS]RE<31O=Q5:KHe_Pd5T9KK?;[<29b1=F+bWdQC+K@R_\/@Z]cd6_+@02fe8S
CYI7AX+Z[aN2ZQ,+IBLAC\,UR57eMFNJD,#)TJ9X.)L,+EFS@B>a)P@BW0TZ[Wd#
ZV)ANY7Z8W04&.JP(GGB;^UAUNgROAP6#>-Ca:4,>f7>,_(b@d41D_O2)e_<2X/4
6R6IU;#a]FXB=)5g8aNG\.+PX=EJ:DM:RVEIE_;3^_IHcG?E=P]5JE9O6,,gGBQ3
BREg[3#bN\g_VT_LSW:[dg]+9^>Re5.E_\M=4(A<CCLKAb,#Z^BCMV&Z@@_2-_[;
IEIMfT)?SEf4;KWS1@_<QK?2g05C2]TLN,CF3Pg8f@@C&;M)0>5B91]8=/b/G:SK
3H\d>G>U,E.ZKH[FB>K1S6f&_1ddA_S<-BS^VbWZdUD->d\:7(D51cNG)[+TTFLP
.eS2#.-RS]&E7@:9>]\dd<TXQ?[18.eNdQc+eEXJJS6>IR4_RN,8.N1F>X+HBVg0
>B1UI/2]B5HcF=EOcS1P1K-B&Ia6H^)T<-0B^[JOZTRL4HICaEI#-faEED+b,([\
R@,d?>TX(,70TP@N>af)eSB?+ed@KefEaON4@WCILeTD0;O?;+S>,XGR0G9d=881
F\,^8L1JZF)8Q.AMaA.:eXJZI3@Y[6(=MgQHPOW)E4[D8NFL>QcT5US&3dWQUd@H
,Rf/NIR,HCAXIgYRI\U_4@&/E#SV9NE(SC:CDQ^gV5=-2/.>TR;aZUT&a#/2-dI+
KX_+<(fIPY(I41LKZHLZZUD2Z<=.RSBfIG+0T>-=&W079S^M6.ga;#;6X:a@G;YY
XCIPL[D4V25f^G2X>-8gIGKU63<4&-HSQWB>KS[YJ_aMOd+27+786RKC&P37V3&6
VW6Lg1FM-dFSLg,+C/=BEC;Q/#VaFB=+-&E&b_/?5#,JQ4JgXLFD-4X9K]\c?P0D
1X?&c\#g6ce\GKE40I<@/6Y?\La:\7)>WPa)I+S/-c#<Q1V:-^f]=g1<-]PP#(BC
U>X^^(gC?1K]S<(5@/2(,H95]WA9(&gKg-E=D(1G@4/aJR4EZZ^-bF6A;3Z+@T2.
PFZJ]_))Jg?f)P205XgT>g2[8b2JJ.5CTQ]b2VZe>8]DSRWH9b+XF]=/7N2VAWCa
\SK&D1Ha>7Hcd4CDM.X@6I_=cHEG5_IVH4GL>?P+U?=.VYG\G<R5H(<W9+bY7E]g
GK\M;R/R<a3<^L15MFEZQ-Y.&5J#c[NQ)I7X9ZUafbU91FT.a3e+Q<aEg_:d_Y/&
0W:P6TU1P^(D5MKDdHU.1cEWOGH\7+6B;ARO;1EG)+e2:aTP7?ON\)WWOPB\:Z,V
#c2]WDf+SS&dOU5^Qae9KYG_AdO@)PHFV+db>Z>?YZRJCV7QIS<f.))3UET1RN.8
HC?#]HM(DS4NBbZ/GB0>QTPFF9]8R:BfQaC)\_8@I\dc]P69Z-V\DN@67Y<&NDg4
;H[Y+3eJ^FJ@&6]PO46JA\3:?.<GV,2_6V65A)_WKT?I](IQMV5e,.]d,d@;aCd3
:a4Q+DfFTZ=EEeT#XeS8+N(f7/Hf^D6_IMM1\IObMTAOF4D58.IF@]W<OZFF2;LM
XE)O/NHf((_;e(:FcY6e--.:BA<7eT0QE9?8L<3V=^4[33UVY^2cg.YD.Qf#9+O1
/UPeQ],30D6bRb=]45:<Q:,M5=&?/QIDJKeF-NG.X.(4:+XGcX>[HD.YY.TKCO@(
dR/9H(2#4=DTMf/;LR9:f;fQZ-fGK2_/KO.9_cgc9EEJ?0:S(L-cR#UO2G>9+YgH
\.N\H(/WT8QTbfZY3(f#P?68,LCU_e=J_?;@+b?^QOU1b=EMI8b2VbgJ.a0L5(ZZ
@1\R>I>#Fg=6--GTK[/-f>#IJ+Z)C?O@VL?L+gK[/H;M\\FMBV?b<:=MQBVGg52B
9MC[B2\)YA^G8<IcBM7\TZ3FKddGYHF&T>1Y9_)]RUBU@O)F^;>[Y#9_.ceYfQ3_
;FcK]NG6aACF45_>CI#[10a^KS:N#57>dH8G.0Z8NfN,S+^c7@BcJ]H6#1&XdIX0
;KXLNW)b[UU35Y^9HOS2/R173aXW#1,CA/KRY2cX;g.AL6342<CIQ@+W7=S^F9#b
BV8,F)<Yge>Y(T]3f<24KDFg6eU/8G4dF/KUb?90F.cE:FXU:;Q<0,e>dYe8&V\_
7M=D,FSeWKIG[ZD(SPYfPIPGW601_0==CdfAcTU2):QC.<Sd=dA5dOKRc-b;YWDa
-2#4aEOTgbcVAA)e\NPKdQJL<RJY0&O0Y&fO2N-T9G\4(8>d2R\3B.STY__Vd4F+
FDSFL9NWMJ(fffWUZZ=GK[^dTe#O&a/aIb?gR,9c2\YL8B5X6^EDJI<>LKeANcFE
Wf3W5<:)IRgaE?D0\A:.9-)L0T6+F;-Ug=I+#d(07H35\-/C>6J\6AQeFY>7[Z])
C[ZHP]@bc)1B,6+@O2d0P8[/S?Sda3=L7/EE9-H?FE;YSSf[VRZM-+XYB6/>KB>c
<c0Oc82d^)-#A1S,>ZQf8;7)BO3,486[TCNA6J[-.)M6WS^;-8_<d)J4971??30>
]M2(G=.&((^_.F9;e1)[9WDXBX1D^,_2AG.&2KFOY+H4#ILIORTV0]TCD+XG4L10
:0EWGEH<X)e7BE93bE@O8N5AaRV[aJF+<fGNFI8M06T<3?WGECT-8FJ8b5YKQ#DN
5HMLMI]>ELgVKb/?##[;cW9[/Ye_fNN\[?[c2T[1IQf<e/4?[N;a9LLbZ_A/(+T<
dN.^JcG^+-V)=23c8E8&9&Y&]T>;4(H(LE5-I6.:6UL;E=.665RYb<aV8<X^WE^B
(&43(8Nb<752:Y)0e1P0M/-QBdg;ITBA-[192FcW4:UI;J5Y-^;:=]_S=Bee@>&_
7@J<&&e.V4T;aDcPGHU9^;DY7C,1)=U&eSY9]1;=+[KR.,1ae9^G>/]&HYKQgYGE
#9;]+Y5UZGcY.,AF0O[d;PI=X7-?6O8H2AgT:P^Gf7Y7X=/a)32@38<22>0XGCf6
3M..=@;--QYCb79c-0cDH8/TZB[I87d8gC:_S]F2-U^N4Qe2DKEPE+._4+Zc@bId
f9X^+T#Ya0/IS^0BgRCJ&:X:QNCIIa_R:K6Ig,_]XPQ2fG<,b^NJgBZ=ZDePZ-51
b1gaag,YKL<3YCY+7]#.3ZQ.+Y:K1\UVD^48Z38QNOI+)@98)6([O49Z^TbR17cA
7H5?J2#B&=DDT)+189&_#,<:A6(eVUCCIf)7c9FM,9O/8S-4Q(BTK0E]DZF4J3&O
P[-e^:=WB]_G^[fO[30P/(O4P)4Pf3fVTWSN,C)e[9AI+)5G^,EMWKT3T]cG<[)Q
L0P:5ZEB8_YYLAA-NZL0CF;AGS7V1cg<0,)6\;?G6bf[QRaOZ?995L3J.VZ?<&Q>
eJKbTQ.JN1^XS(a_Q[HXOME.bF]4>Ge.NL9dP>]PWIOSO+OW5]M&W[IPEM=Z]]g<
Qb(aW<X(FQ_&,V:fDZddN@9L?YML>-(?ZYL[eA+QPU?g&H>(67RJb[?>[9>XR(3W
@8&5\?1?V;&K@0Z_P/G5#/a-,ed4@0ON]=X/2X<^^IB9MBTc,f3#^gb#DAU.H_0B
D<IL+@8d1d5QDE)5aUS\L9a6)eHL\;:9H].9X\=+IeLD>.O0P5@c@X6K_EbC2^Bd
).85R]d/ZTEDM/;ePBM2-X1Q37_UAS3.I,b\@g]XSa0X;f+E#4aG:ZCTHGgP]_&3
f6[PDgL@d[RX20:PM(5IIdGg?\M.g@:QaHaf=&^P)<FGV,.&9V798Sbf30GdN4GE
O\=P\2G7gE8BK0]dSe?OIC\BGWbL_3:&LOJ>3a5?K)W>b>H/I0U.<?=7/D#(GbE]
<<QT;X1#PZQH18Rg&9&EM0M@V@VWEQ4,P#?P<0(_NOSLc5.CD204OJ>IAN[3NaS,
L7I9Y3W.7;NYT@:AL&G/CM/N7[TT,g#F>C+?YR,WV;ORP16+bER62I43Y/5RY0EF
fD\Q^&fBaN0I8XBgW8b9E+D-403U,gC?_<WAB<.Ra9GI0c6gD4K;E57RDR\dSHQa
Ue_N:]T=3K67N\g>AR?;>(N;W:KAX1K:1EeM)I5g2@VbJ@/2131Da(G;fV>g9Q#S
77EW[94+C>6^24&O1U0?OORKF+BYNV@<REg#2WNC]L/Ig8KUZfJ-bcb/VS)0]E8_
S,;IB<4,\P<\cH2N2)b=cdI;d6X8.OXB;M;E>N7.])?8G7gC+VTQ+Z@eKOIK]E]8
+WN1+8]CbTdI6/.XN?aaE6JWXK258B=SY4Sa@?aP]E8,ZH;0A_LKa0ZR6c#Y:_Z-
O]Cf=Uf\4RF23L8g.bO_MVM9H0YcTXB&#WYP/:aCBI,+5[]Z:](]IZ?@?dEW@>J-
Tfa;OU20J8X#Nd.FD8dX)+N;>2,#SN,UaKBd-_;F.SH+F$
`endprotected
endmodule