`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 1000
`define LAT_MIN 100
`endif

module pseudo_DRAM_data#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/DRAM_data.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency, 
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:4*64*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 1, DRAM_W_LAT =1, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8191];   // addr from 00000000 to 000203FF

`protected
d1IZY]/65)^T;>gERNX^;Y>4(G@f,WJG?_bL6e0]G[8UA1AZb[+T/)-ED=R5,3CK
A@1.[<6g^94BHF+8\JA(8=W)Y1d&a(I([1.:1PH3--([7>]0@;NScN00?b]0ZbgA
dK71#gITKN??BYAc]6[=Q74SXJFgV&HUP2\OWF^S2CHG8&FCFYL/fg^NUVC7ZRN@
GHUYL26ND7Tg]]Q<X7gQ;;E9@1JOIZ(Ig->?3I+5+I:R_cW1LL?V2]d<&7e-J-gQ
KA(297UAgCTTD46N-R-666Gb+P6OQF4=LY+>\)5R^YV:.6<0I@g70UH5X2ecQ0^e
[/,d:5=SdW3LY:]9OHF[e(\-YS2Z:)@[7\;9+2@/3L&Tb#QXT7R(e_Z4c+5c\O46
aLLTA83N@8I+8S+>1IQ3C?#4I)^GKAIZ5OBfQ\;Kf]6VYfDN1<N?EN>P&1S^M,cZ
PdSZ9IQR68PTI(FfPA1)JC4gc)U[=TDPBEKR)dNRJA7[#Qg?ZYRd?D;Z-1BZL#W.
\,6L8I\D7F9NU@UCYB#9Z6(Q2]GBeN5Ne&-.M]413.5PA/eAcZ.GO0.<Pd;[W1(N
T<;<E]L;R]4:N9E7;fZ<H^F.U^A@6g0J]8;(1Q</POOJAQ;,_1JD4EeK0HYJN(RE
3^+0Z;Y,1Pf0e>DL2OUJRegG)&O^=51/3[3;ACQC9f;>CHBP@D@/84Sce=4#R47-
EZ/H=:;K6W>af)OZ3B]dES9>X:d5I:7=;3Y3Y4dI.L\&:]&Z-/P_<:0MTQR\U#L;
d>#+9Bb?+T[/Y@18U^-==UPG_g);.7OH@2CH&<02MZ3c:VO9>V2X(.;TLHG=He-\
b-XUaIZNRCUA8)-INLECR:4;@0UW9@]]?ORE8<AA@Z/7_V8>:+O,b;=Q2VJ<[K^d
0Z<C)>[DH^L5MU]QCC@_:U[K.eZg&\_GLN,=cD6:/cYL.MF#0\UfaBT&=d/.:QRC
52?Vd4Cc]Zg?KFV/b/U=eTG#a#LfRg.Z)-:;c\;]ME3V:0f<bKN>f8PBJ[=F2_fD
A/4PccV-@>5BP4F;OQ.-TgaG_OKX6&fYdeW4YB<g\\B@Gc<B6b#O1JYgc-G^EQCA
<@I3cV>0/Q7(5S0dKR^;HJJJX6;K&(^JL?>F8&A5AV?X\5#2H191XL_#SD+E0J[;
=+XUYFQ)c^T7P812eFBD@dMB>9K.J21WQ>CdQ7+\f@LEGb&c>=WgIQSQH4Cf;fa1
\,(AK?G,&f0XKb.Z\@<M>SQ5QdKH5P6Q.C0bAbGS8L4Qb^QZ[LG8Q_3K9MV/RL;g
YL<0,_;Q,?,O;1X6.JIJ5.&e\aNXHO7E#2MG4GRAbd))4^O=8S7S+JMSJ\Ye^LD(
/WaW1gUI9H[XU6b:G<b8#VV8NJSbD2eV6L:H77;bW3dT8H6^7COH+)edbT-;S3?O
b]G>7CK;V4d>(Z]@Sca1,A<O[e+<AD<^2E^I@,^e2YK448^I[4GQCSWH/T?<T<LN
KKGBde?.V6BGTI.TG[-UcTbcGW(?ND;]2]Ug5C-gD-G3JQRG@&9CD6)C:0V:>]gW
=Jg.-/1E<<DPB.E?A]QVDM980DKZ11/9STKBdG9K7H1]=dAP6#B&D5.80R(aHDK?
f6^SIe]]^LH1=+DA8I1D_aZ5UE3Ra@ST\T]B)[c)2;SdRb]cR9&40d4U:a)H[#[T
eWgbEeA0e+:cYO>XW8c,1+0g012FB8;BMMM_/MXX#9ECSeAXJB8??bT=be/=.A51
3&ER_e?\,d&5(+1H(D]-AP\AQbINDb8[a[9])f-,H;HEZe7#e6]Y57#&E><;;gb9
>2OWA>2HW/a=UA-ITGVB,C8)bPd\aK<].ASBW(dU=/^:bVA5&ZN\QgEJC5gJWFPK
<=<-1=Z<a6T2S.SS;=PN-,Y(R@FWS>:1/L(9H55ee<UT,K?+a]UE:d6QbeaABD,3
&)18-DTW>2BdN<\9?e,U>X@Q./8/^CUH/SD6c46>>e3)5IVf1>RGB-&7)K<b[UZC
B9OD33GEDOaPP+Hd2>]7T:WC=ZOSDZ@c[e_JSLUb.41N:8G_?d2<#P]^;O5=72df
f.00FQ25&g]]^ZT,bJJDD<)AF)E#_YV0HREJO/WcIZ?1bOGI;^P,3b/dE:(#S9?c
QWG;+//c)g4Da-7=@N05W+/(JLYN;;WHC;5FU,@M8,2b:bEA,]_6PGac45HPMO7S
)2X]a06S+@gRUg5@R&0c0(]I84-JfQ-;7.TBc]LAI]1-9749E9+..XDL=^;LF;#H
E1WfU:WA[54U\4Lb79.deEYPACC185)<7>NO@J&B7P:DaJ6,7Be\3@+:2a1#_STZ
9=GLUZ2X<;GQaA0Z>:OPR@H=7EP+^L2_YA3eV5^<VV]g#6Bg#DV/cD7HdEJ14-SN
#,_ff<^bg9aRbFX+#2OOdM:.aA46]d0LQJ-.A,Pa\9/RS,62T5LEWWQ185IL3:a<
N2/EPaYP25/38+TQMN3,]5GCZ=BW>c(CZ6;,46_1T:ROJYDJ&c.<e,P/FaEaNTE=
EV96MJ/X?+aF2&92IS5AU2@N5?<1\.bC-[.=ZfI\=LI?WYYN=W3G/eLUOef[U;/7
LI+H_A(;cSR2<#8E=2:#-C]S\S?8RRXUB(7O[cBH0\&EB(\9A\^9T.[=92CV<+8B
ME,gATC]XZ&->M?I#_F2La7KL=YO83\Ubc?>&,Fe6W:L_23F,X(UQ:<CH/#PA7NQ
C342[6DFM3=,dZ>TMGcTb2\gZ6D<=HMR_@?S<-UWS^A:BN0a4BRTS)W/6A&C.d<O
;:+F4<#e>(<JPK6]<_PCbU.(CI4Me;YIHJGM)dWMTO].,=YVL;1B?H0FLV@I^beG
JYcf+Mb7KEUWEH8/RS4-T]54][8VFgGKFEW<]BEZ#K=N_UFAXC3aF-=XAG;#LJDD
J0S.?AYYJg0PMAa500RENK:LQYcRQ2W9e2C&=TKbK&3-(XCS-QSAF1LXFXS\OZ(O
F+P;fA+40a,6d)768C>WPe8DTVC&#0I&@&g)HH_RB/[QU092:56]=e[6dI(D),>O
1TeeMXXNET9D/U.gH)gRaOc/((RdP,99NSf4WRA])gN>HDKN6fLD1-VGe-UYaIV2
)S1Qf-NION2)NHYX^8T&T#WAP62Fb[_)YdW=ad?V(2PCRBDAMEUC>2Ic8Q=f&/9:
W>Z)O0Gf^\Z?_PD8#_GBU@8)6>7G4RGbCa3PcO,QJ]bLTY>@cgJO,3]3(fAgRU2,
8T^3:?S#-Q7L[S]#6:JZeIA#D]f0)],,WF=(aE)PVV^]ePa.a&fECA3MNXaJW?AH
SEeJZ7cMdT.UeY4JD80]ALc/6\Gd3;I@@LRe2<3<-#U.5f1BCY1W16WFT>M\MX?;
__NW/7bDYd3@Z8QUH[2,W<bJ4b)gGTaaI(Z=@4ee-_WN91?&P>(NYG[6O,f#.R@0
H8ZJSEBL3W(O=+[CNPU-AaR9fA9U(A_WZM=>(TR11KLbRFR[2dGM3_PM[PFHO,K#
@Cb;MSJ38d&&&;WgH@fS9AU5dKE@UJZAVQ+3Z=)W]>2Y8:=;V_.PGbUQcQLMC=Nf
;3K=&7aV0C0]?CKO3U45./UDYQV1>0QY1Z1G6;eT_Xe-.5ZE74a\HcBZ)U-Q+g3-
KS0Y4Z.205,-KN4-.c:;YW/>LXU^C9V6EHQW9MN:g1FO_(Y]@+9[J?-&b,&cY5AS
,B\E2E6>:7gM(:X3JY+f\F9>d4;1D4+=K=>+T)W,/B_#Tce7H0aGS?M2X@9=BQBd
V0JH@E=>TFb6cf.9IC,+-,.8L<DNAT18eC@;VD-W=/e0=X:4VP7NT5fMH7A/.6@c
_7I_ML:FI;];A1@/PH92V=8FWbDARUIB55&f.Ae@CZdZ;\,>?gT0;eLda&K,8^(g
J3ET[d^_X]DCaR\DcYa>4Q1fY,7RTGJG/aCB?9(,-[3ARDGXGGZbH<T)39^WS:3_
[2G;LgRTL+,_e@>e:de.0g(>#((U0P)#5B2&TZd+0Q&L4d=a_OQ]3e5&TbTSYAA?
_F]V)@3@dW,RUX91IL,X>e_]NHbOZ1+>51(&7UX;2[/1#0>)7B;/BP31b[E1SC3C
,^Y.dN7;RKJLd-0/LU\]SHF<95H7BOQI5&,,<<:TVWYb&c2MY)#SeIX.MKG]_Y_4
bPJZDd]TPH<JC0OS0<UZZ<[+]0AI51@):,SgaM[^WL=U6MAd\^2<d;8)SD)_(3cE
ETQ]B2aVF=C&(baJ\O?=gYc6/O/g#,>gCOCN<a\@_E9?0ZX=30MgM<@:KI5-X76U
X7^_EfD1(?KQ(5YFT=@/+BD.;UR1>[-,,P3/[(XUba?UZJY4Q1CE.EPH,C;cLfdO
S>UU^L^;S53.<e#/^^)2]]NeR)JBUg5X-8=gF=\M)J7(P3SLB@<cZ+6Y7,.G)-Za
E?IG[(8+bP4d5B6Y/NfRMGNA:a/ASDAY&f]<C#L996G4YeW_N5O#0e9N9(HZ[-3,
fW\@PZABX.Mb/U2][DRBLRJ6E<g_UMA>7ES@)-8gRL=d3YEI-d^5PIg]Xb,;.G]H
]^SJ)fGUW]->b1<?+6(82a)1e4G=8>+GW7<bM@53aUX0,ePW9))E)IAUU2Ke5^>H
X6;8NW)H,8C_Y&_[/OQHXQYIJ,8H?A0(ZLM)U@Z+DdKLS-O+AP;IXF]084=U>+5-
\?::N9-Q,IS-&<U@>g)Y:OGSb]1Z4;4O<Ve-aSAF6bc_B-+GJ=Jd4D#D/0-NPY=:
FEcJK#Y>+#[[WG?5f@9.A_;DX>gJKR@&RcL4<-)8A<SH5?cV^a?<_V^(HHT4W]<d
1=67F0^TK:2D106MQ9T1W@\5/LI6P-=#96f-M4HcZK[TB?7eSKa/<>;bM:dM0KOE
gHVFVRWaXd#?U@AaW,=bX-SU6Y-fD:W2012_WLF#?2P399/D,g9?WMe)0gcZ^K.L
BJ9JC.abPOGeF[Q[,V?^#F>NLK_S=BDf7N@AW,@X.1[0BJ0@.HO=8(#L=/R9Q#]]
D_X3?K/XCEe\(ANR&;SY]J6P;;GcFJQ^<<G](;DWEb-D63(fPJgV=V?EIZ[@Y+D&
OJaBK<fc;ODD6Z]c@Y3=8J/]>D/)/42d7?]ZAdW+f>OT^A6#R?27_PQNDJ>.UF_D
SP7>TAY<HIT(A<dJ3-MCW-:-673XI1FKNW9//,;^+7Q(RgOc1EIN6-IW&cL<O@]K
)DI@9Y>Dc]T&JLVXFHEda48PF\L[IDY9#e.S+&B2A;&A\EXN^&1WOE0E=64E_F[^
IdE-O[8ZJ7]f4,)U:TUEK]-7>0^c3_?T>7@KVJ./D+9\+<#7bCgVCdP)@7SMSHJ?
@4H0d3\BFDNL-F@0UEI[>>,,V1)I[LHSS99^+e^I_#39VZ+H@/=E0Vg_g<0U]V;\
/T,36-YN65;^G@63QGXY?@#8F4H;0>)8UR,e&\.JaSA;Xf([&/=@[E:Ug7bB9GER
C7DaMg#)S#Hb/#V,GdL)d]2U\WUOM,7/W7=].9d:CfP^)+d1<M&.KJS@<^6TF@QS
.ReS1>Z2HPJOg=@A,N@1N?dd^7?BL[RZI]9QCA2V@(a=7dGd7E^Ra3@NGGgO>_1Y
4/++]c#.55ZYgZL.I=96JU4.>DK6eW-/G-L):C/IJNVF]<;#=ALXO0,^7>\<W-HU
^O&f1d?BC9,#bQ.WDQ[1]_Bg_Q9NgFb/4aB9M8eYT562F;]gD:-1]-E_W_-CZEFF
LQ6<H<RU6F.K2<cMd^cRM8O6^[L.PTTaAX8B6Ga96YD(b0H64C>Q5HAZ5+,VHAIB
_32V=SG8X43]#^f8aD-;cXYM=G7H6cWDc^;V<b.:8)B/Y;:;60NE\7+bagAPD;Mg
H&N8&&H7]]8]Rd\]52VKMaH=6)K+RIF4V#/@+QV4S(B.<0\QB0CV\R>+AG#;4Ocf
]31/>7BEB3<V2;cOe2(O<[G4YXH3:P.E&FUAJL3+I[[eUgY-N0R->B6Y?dcRN,B8
H)a6D#RCaLHF4;7IG=VL.b[+)^I=aGV:IY/FT=[XSW5ZT7>cGD,4Qd];FXYa.\F&
.UYed-8/A#L49DB^(CNOEVRQ/ZPR:b:A[8^8<F,JWZF^g]?(>F>SOM5GJ6VXAF._
d?_H4@_a]X]-R=C&5+6F.P\0WKWLYHM;G20-+(;23<6e?S5GSKQf6C42N?889@?_
86TeU.?VSEG0Qe2GC3e6^<1@Bg<I:5[Z#LAN8YNc;BP0YL#O)VXXK@PH#;NJ)3@&
PM[VNEOQ](EZW8I0L2b&-F)^@Pc=_NP/&f3FGf2U/BDH2(,N2&)fCVULaN&,A]]T
)15IPUL<Z\bCPUEK#(ZT^.P)XE<;ILQ9UVJ/=3KBYb+\@F@S-/<O[ED7-8Z?>@dK
?^3L@.W7BKg@L8fS&aP,:2G5^LGGES_;g6,LMU8),EUI0SH?U-H9,4K[#(cf6/NI
).;+824>9/P.?L]YYLZ?_S=ecHd?)WC]?abRY@,?47&\Y4<+MVBO.D>E,UGUT)J7
YN0^7UTF?+4W\@T1?5-+VNTDP>Q?\d&\9STg?PW2cWO40GI:W)V?93S@6QW8&0YX
g_GgRc4QB=f&9T)Q+d3\GJ>&.F:@;2WRE6.1&>\/cA;AQWNK6Y)R4\<F.JgEG_D1
<O=7-6Ff)8+LL.N05-ZOR?M1Pd_?gEL;.(TU>32NNdcFdc:BV87dc[>:7PYOSL-H
>EU>DSBDOYM3c\K2E.<?8YSROF)UFVIX,ZEcDD]Yb31J8AI[B^3/PD[_&M>./OT,
B+],[0Z)1EVH[b2^+OCKNO#YAT4(&8/=KXDC&)8eV#c,b9fH[A#e<#,_F?8:6^KK
29Y(JUd04f?N2&QI=V/VJTY\aCe.eV?c?97_M,CCFFCVVYMN<UEPO\:KZT)NWPcR
KMMgI)H9RfKg44#X-b9E<f+ZRZf47c;7YLZ]JWfNd?-)[R[/1d,.c=_Hag-[)=FX
9-/g\,QQ^X3ecRNFY<JA#O]eQf>g)=gKA573TgX/P6^U8KAID\MGX@aRZGL_8BI,
.#HaM[H1U<968,b/V6?,/V<NJ7[9XNFD3_D6dXf,=8K0+\VR:6B)Y-/:@3YHNS=T
]C7?B\82Ub&V/WbM@Q[b+U2McIg5[B0^FEPHA/-4UgYG]EYFZWf4LGGC<;-N&cdR
XgR]=5UcM<9[?FdGI(H?I\eC9gKf:b^-GKE@KAG?.fI<Q)MYEQC#/]-CS\DG6MQd
HGN.D<FY@;HFd\.ad^GUJ8YUC6SU>,:OUgfPBLc&C_:XA73Ua+EETJK3)=--8bN3
]ZY)\]9Q/bW7^CbOf)^5M9-:@O;=NNG<)<Z2cI\TH:AdR):WB86@YC;:(^]N9<C+
#XD/<2aC]=T>SaTV\aC_3-)EOA-W9B3+<8X(S:bT+?0\d8XN8?/T@R(>LIYCI2NY
Kg^AFS<cHGQG9#5K=80b-O,95M((MRf77:-eNMfKfAJUEMRbg1VEe1cG=0-+KT.\
I5&1J8?f?X^Va<>5Ng;Y]XXHa)598XcVHO#JdX9))VZ_WbZb5g>R/0A(TXQ_HF&^
7@Y)&#&6\.:3WMMG#W+WedGQ@20Z8ES9I.;3;8b2^3&,P<85ZL6FA1Y]gI7N;53e
;>)P3RTa;d1<?-535a\D.F&9Fg)S+O[6.0ED5;d0->+d7&;TXRAgXWcV7Y:K:O5+
JYP0?BF4;J17.,B0f:GJQ1<BfM[SKa+A>0TJ)DT&D]a<(.FRZGFV2@OcX^TG91R>
@HFZFC_\5?W6Y>Pf-;8ZE3e/P2K6FNX8e04EKEE6\@7+HN5bIdd<8fM;d1?YRcg.
XDQc)dX(1<?#N1E6_+BX]g)<\S_DIdPV(::O+Cg,I(;dYYc=gYSM7fO@3>[,[Z78
/#J32JbQ)B]a?Y_AF(=0OQG+/GOABI2RcE)>IY2T/??QdC3YG)dT>?,XeC+>EUCX
@3N4#g,AHP81?eXW\5K(NC@g>I3#>)\,=N8eg[DE63C>[4+7DM8AfIXE:ULA]1/,
Wa,Tf]LCT]Zg-+X@N-UdaCb>/D040<8fX^MCZ,XU:,1e?HL(>[>UW2.[d)4NZJM;
Y=Y_<XM;374,J?R27V4c\5?fIKOI<c?;E@S/,0M=QCML[SHae&<.JfB8a,3fJVM0
M3GM[D#1g_b\I6dFM71];eND8QbA29(UBJ==&,H#+ZaIAS-#db1OL#<dD:KL?T3Y
g7/OJ2N&FWNC]OgF>>L7>;(SFRWU(ZBTee8A4V(2SF,W5106K)U.6<.=0O&b.;L5
>APJ,FbgJ_(VG[4Z-J6Y\>QeOe#eR4H3-TD/@>6-e_Y&A>#f]EOQc7:#9LW&KATS
e?EL,=bI+R;CS0:U;Jeg/PdO5?BLA@QX+PbaZ=XFe,OILHTZ7S2-a]<5DSPNgVH@
=CG4Z0/2S\[2&&HTHQ1caD_ccEIB_:g+(A;RGL2b=XX]>4Ya;BQQc),LJM,)4DO6
Yb)YP3P.P[aD.\\0(_.HU9OGYQ;b-WE<LU8;7XQG7IYa/1BLdc\5bg9P1cSZQQ?3
b9(5aQ)\6g1C&^a[^IW:,UE>gJ\N2fL=JfeM#&J49NT3[8/5DQU=Q/cU3#KO77:/
e=/#/#WAbBb<2N7K??>KQDM7H)?S\P8U&-If8VXLU]3M=#EE+<,^3^I+/-MKL>_P
CW?gFUQ<PE(Nb?KA./#7OF&@4XKa4JdV.<K1^VI3LL;3b+a_S1[NNJ?,KVLH/RVg
)Vdd,EV9:?e(Z50T<c?1,2NDBZYP93KC<)#\SCGS6[?M#T8@N/V[g884d+X\#_21
UZMJ;_a:#_NWVaNL/&2(U<-1IT4RO>,\G&PQa?[8#A-J#E.BJC1.;K1CTQbe&203
X6@3=[_eKaJVG2dQ)^@X977UW.U.<159:^gME@B8;4NVF)EHMaOTLd0a_H_7d,J(
d9R[AK5VA-GRIa,>Jf-9/PcTL1U4eAE,:&0@276KLe#]7]OeB9DI-94H-ZPZRWM8
D<afXKR[X#LRD?-?-EcUOE@MA)=<<:/[.,>EXT/=V,@GPYbUV@17Z:W#_IOM\Q/0
H&RCVI+B429d@4f,4b/bgGWVE4OD=Kb2Dg7JRd)49c:J=]Xe=F/ZfRg-TYO-/258
bHUP)U-K?3]U3[FI?KEAB@YYU4)=._=]2&]2FWd1OG&3a3,@@cN,@<e27dH2eO(Q
3\5<c=-\RL8A.@P)@E.dWG1]C-Y@E1Ac&C>H^-PI2W<43LAQTK1a:/[eEW1^W6KZ
HL\TY81(.Wf#J0O=>V=S__0<I,Z<K[:4:6D6LB@X,,b008fH\LVg<>:[bf[C-U12
3;OCZdaX;a33?Ab(EcMDd@D7X:eJN_07GYc>X33@5c;?f4]2a6(X.E&(/?8dVf90
L#]LI]e@,cEaKX6;K6M<PgO/bZI<BMT6TEBIUWD9AUf;5M<BP@KG#YO/;F_#I&:a
_7-GR9>XfCVg65WGUdVO(9fDGOFbEKN6QJ&f3G=9.^VRJYM\ABN)KA16:A[V<bf6
GfE1^W#bMJ1Ba7?;QN7,,0YR_CEH)Q>L47Z5VZJ7UICMOFD:NG6805(1PH@.ZUU1
L:+:NB-88S5b0CaWe@aN9L^RCd/]G4.>#5E#Z8^;I#.4(NJDcBQ_D>5d>,SS0,@B
^UWM\0&Y2)ICfI2F@+UKa),-.Fed.aVS7Y_MdHE5\R0GJ<DGKbQ#O.OScg5(OGL9
#W=@M+71bg.;88H?KH-dg/D8C?0QH&2Y0R78fV&?gA7f1APA\fW^FT^6#^e3L+Q/
S_5FMUPG37\S.YN#B8[G?)1NL[&B7P=-f6IDRb_5#=.Q^/>c89?XE>1B?N#7Jb0L
<4XL(69,34:+N4<9\540f@,L#-JN[fbNa-A)RMN<1:KaD2DR1)^IEF)L)&RLD/7=
bG0#-IC)0VTV_Hb8)O7D&2NG[C645bLc[ZJ.@eIJA?K8_.^>ZTaMFPC#-2;6d4W@
>U[Z-A&ebTO=9+WZ[,V?/8BaX7AAF/a7WbT(@M5I9DRL5e(VNFI0_BdC3>5V2ADK
6<F?)Rf/Ug9&.PLf/0ae?M=/aQ-1>A\#OfW-8E8R[62gAN&^R>E5@(:?+F@8Jd]J
K:L=\Hd8eJ>[+RH0^RHDD,TY:\G_#/YJHME29U/),2J_W>.4)Zgdd&BC=d\;@<CT
TX99@-_>GgQP/0+N<+aF;WVD/I+M97COG57RF3\7^WHa]_U?aMYb>LD-P^87.@\D
=S73C;X9^P2.Q<-)TPHa\aO75>L<CI,Ad>Z24;C#_H-0a=1UG:H)MG#K;d7#I0>8
<V:=/c?>\?P_RWII</6bAa@V0_7Ie5a@Mc:g#HZD,_Y/92?&,^F\-J^#bbAN\YR6
(IIQ+&61A./J76<9;+UW@6(B)dN#d,EeLR&6?4+;LF#NK\B#QS.g74c_6\NQ+_O8
f@=S0474.[f7B@5FNdgccDQDVMC800U5E4/RBECcZEa[YK@b:4BWJ@Me:;)c-]]F
>NSQ=<(DW,(A2bT;e<2/FRYH5T6H@O2N8O,D<bOBbTDR5XQEWS,\CRgF-.5MVC1H
^TVV=D6&9_VU4;EL_<^5/#[\+JY3^K\:])C#0)2=RN0DSE-(PJH1.0K6cdL#.e;/
W9\(+TGd6R)V9Fc2fE8a@Db3?5a>-0\B4K,McMe;I\Fb3E<YVE55I=2)/983?ga4
D4?&fFZd#cV,=HAVg#U5?0L_NN;XBA6BQRA6T?53UL6d42QSTHcCN<N8A[U[gg3&
&A(g-cGfCQ+?2Q;+#/=NIAZN?T\T0&<,)DHN>SN\eY?ZJ>-gWTN(d,SPK>S87J-b
:X\E@..O.eB[3g3:2[H=BK5\)a>@-?=]-eG>SWW?T#JMA)>GSW)Cb:/7PHHbce3_
]_gF?C@@g^FHdRaGLCL&+Y[U\]K7#22fCBB0MK3fH;VP72(&<<\gRe)d0KYNBQ4c
MgJ\E@.dHG[g]L#WA7+4W81B+]Cb.?:5D@9C96<0PgeF7dB\c?/Dc;-D6-CJ)Zd0
]gcF=R[[<6.H9.6<6dF:Z^NB;TFf+?HN-GgUc8H4NXQC?0aV8F(B_F?_.\:07D)[
J&WL_=E3?BegI@+G>=8497a8#[9NL/3A/&JN:SATg#I\@6,T=3=P^RA:[cT/X@U&
F\@:YNTgUD:?R.2667&/ab#5H[71>[^4OK8RQ-fTK-#@XD>E\(>_)SbQL9]Z\XN#
JJ#Yf<#A]3W:>e=Z:48O.UEgD6XYKFR0O^gQ1_;&dHWI-N?+VDJ,OKd)-:R;<f-f
.IZE0T9&M<X]K6]C@_7@&S..#CZ,P[e0\,G].^F9ME:Te<dN6C#;=?0ALOL<Nd]]
)GOSgZ6&M&C]4UVZ]b79U1^JS45@#??S9Ef5b^IM0TLJ)2--9ZLRe3O+^&1Y)TC[
25,Y,@?0NKXSVQE2,IG;:@QSIL5I.dg)DX4[M?==J_:.?dAVXJg2H.?bQF==f\df
6^960_3?GG(bAU^T-=-X=5/VSI7+YR[RKRJ3+W5R2a.Z(f?1T1H/K6^^T_Td)S[V
MW7^?\&]^(Xb,UVV2G.,c<Od[aIf4<4\TfSeC]2<6afM=FeIf-CeB52R952N-G<E
=E\/@5ccZaYW92M(#D[:,S_)/6LJ9XF.)29HZTUb31TOVK3E(cLeJca7.;T]8Y9?
LSM;?_TYINgH;?0RTXca3GQ1<1^&)])1SYW)>E4@;6(<g+e8eH:c3?G+08E0VYgX
D(HM0EBTR)6X]Z,I58?YR=V/KF_EH)V>dfL/]A?6d,W<gZ5&K0_/&?8GBUKBKZ;g
[a])_Q-J2P5AFdGCaR+LKYZNF7Y6fYb?(3U_P&aZ913MVA?R#2,SKg--bC/II#N3
)WDO?,Q735,_fVa5>@S#:Le_.b0]@>O]gOe==@(8D?8LO\5Zc3_\=BHCb>URYKee
e<c4\<LO)e\<1<=6<EU/[SU-5,?,[F3a=ZPXWCF9_Id[=;8FX:=<=eQ_4IcL1Nd#
0R4-D@L^?EMCd.&;Q50fQ/R^e1N5e.T+&2XdV3SO146d3<F\?=STg2V-ATS))3CJ
3aDU6f10YK:@e52Q:34Lg&I9b;^WdWb&.>CL>&Q#+2&9>QXE>g)ZM=_>-\f)E?HW
LCb(@]RQT3+X6NCW7JH&N\XQGP86F\KNf]@b67;CI;UbCG=C>)Z-BK#CcO2CA/\)
A+afRTDKQII;+>=YWD:BRbca[8=e=d6H&0&ZDJ43(Re8R/E126/J-SI20JU9U-A4
9GI+VX<@]K2XJT0V?VMg3);a-(L](d_6561/;K_HNO;)MAd142T>aFGAc;0(,N4V
XXEbZJP:[OVe&2[>6YKd(ZYaG9d3PJ^PR[D#;44PC;OgS;Z04N,-<fVg=--\O9B<
H>2J2>0#Ef+?QbUXQQKd/g3aA4E#916@63X2,<O:60L-T#Ee.54We]K4F]4?ME\(
[E_]WZPSROH4WRNNJ].]([[AW3]d)Ld4NDO?0dKW?eR.;_(0@(PWa_YfJDF5)3^<
O<(GCUE?@gX(a+TG8J4ZRB&<R81CT(&(E;3b;K&(F)4ZCE/_d_9cI>U=PaNdU0&_
05=.Q0D\1gCgXN20/g,U).4Jf7EZI>7cDLDU5N3M+A<GWFGAE]-38G8DB7-@Q-Td
EVfXG)85V:6X-_5QGW-7ZadL3f=O(G2a#@WN;Ne#WETMX.7NA6[93&I)/R@&JU1R
CD8c+7cUIRb-5GM4-;d+N=&I+9d;G<N);W@>A;AfMeAT]_F_I&Y?8X7:g\c)0da1
0KPGLeI,aSS+=:^PKR^Tc?.1O]R\7(&(=O80D\E9BPO9BS@.6DBfFgMC+b2f>52a
OW62FB/WR)fZ#E(;05&bC:<:3C)UYTH^2H(Z;(cL&,O@(+UT+UZK]P63&<FTA=K3
8EFc4<H(#dTMaGV25^fF;LHB?)7#BME?X/C[_0.d8O3JC4XJ>cQW-02U3+&Wc<M\
L^-^SZ_2[]MYIC/#.C0AVP^@EfCD;T8e:J9Z5J4YU[,F;3Gb2=][:CV@Uad#H)MR
]9W;)cRI6R@8f@08>#f.?3/8Z,SE<6DO6F@6&1EGEQAZO^4P@1&]IUY1SP?3eLHe
47Y;cK0_1\g>(JcYTb.]d(05C0P35.&S.g[e6JNF]Yg,KZL?^DV\)##[H-<:CTe5
9De/#fA3_(H7C<F-W5aF_4;U3>\_WNZ]BVH,:ECI/GW,a]4GW5aWGPaMAQ<#T.HX
1VgJg?4(O)Lbc)E8;cbc(DcCW[87@[4)dQA>CP/QF(D5W6gc-f6:#N[TMLW@\Y3-
(F0;(0bgA[.[+3,BL,UO\c3G@3,S@-J#^\9YR>)[T@EYQXVbRea]07X7MeVF8D6)
U+\5a;HD:H[WF3L=A-]GGbF:;MK9CF28?1:JV[VHFcN,A:BW&+dF,V]Ke78SE<?6
E[K[M)<HaH15D2^+&@Hd.bc<Dba7L=5SYF;14e8RE]YC)2K\6d@fZR-f]@Z0F:=8
>A6.U2]6<gKVXe+6]f]>4^QbAN6VN5=2[P@ed^IPR[e2,ZI_DDWSM/:\MDea+7MM
+[XRE^KWJM&AH\0)&9OPg?./cO2O)+X?N]@:<VZSK2=W2VG)5.V[VVKHI^EIZ4?P
^V_[QQ^.-0>D(1EM1DG,gIP1OSeI&JWQ<G:HBFW<@Q:9..HILDE<;0g)LfKO(0_E
XO2BNOO/XA<fA;<#.McKPG5/?J6?,VQ87WbgWH8XE8U]4.K2TS0\KJc6U=ZOTd,:
DGQ6^eG3gAAe.:U1@#E.X;,YVX+.7R(;X8a90=8+M,R>Q]6?>MM(EQDHf(5.g_[f
1SHeTI6CWcHZ</PZ\JAU?3J1A^M:])D\DNKeg:b\^:dK9^,9Y(1#++3.YQ)H@;#-
84cOgY/1/Ke>?1[3UT;C6D;KbL7dc[1.N;5Q(EIcfRQ7K?/)ZD83<V;9P1f[LX@W
1O[\4UD3\K6Z:>fMc\)0OV3Y#S2IMGL55&=(D0@4Z/DeW()IZPQ0J9G&X7d4&0N?
<H/f#=P,R25=/L[4S]7\^S_OBBH&/R/N,?;U)0S9AAfQ\d3IEAXcH^@O,C_H>OCN
NO7&YQVES+Z^DT>2F:-4O&f9)[MH_1;,1I2b7bD2WG)]IL9M,e32PT)^4cAV^BRC
FfYBA/(FD\gUYAKcaZ00^.E4\/^XQfY5-b9PPXed3>YZ=5(AdUB#E8(,65-+6KM)
W28#\3&YN58^L217]IBZQ&KPH6(CU&2bLQ=N]d;Z#8Yd2P9+5377U_WBc^/&Xg4[
+bZQa]#F>EE.;<G^KZ_XHDY)P,6LI-S^B_)=S:VIC+Q.],5f>@cIcW-YY,=-cg6K
RG6RV=(,F@K#]<T;&8cC3H)RWR70N<:Yb^0U@9QE#LKZ-4ZBGZb[\Hb7<3L9^>:#
4^aM?\D&SbY#O#1:W=ZH)2(B,#P81?PZPa\R;bI)#YWg+D,6&C5PX)gNV4QMJ86P
090g7Q]YVPeND670PP74GS0G?JBc6I=RD^LVXJ9c&-K:cOJc8Y?Y&Y0-PZ-A_bTL
,E^FVG90D>A8c7_^R1U]Q6f\3]XI&),9<AKa1fV)BM<^V[&V(RYMB4P9H77(QV34
Le-28XR&(6S7>NI99:F(4YBG-,g3ab:.D:3)IBGfeGGF9NYN?1PKFLWaAIb@N1]X
F0+^KdZef-0c/XU_:eP2R9C8Ic)VQ>&8(78d-9AKS=7-Z@]QMe+8g6b6)+:U7Og,
b96:>Y27&&b>9#D_7edU)B5]34<<?0J4]A;]IIHSIU/<7O]:@[A?,=NRA=[QQS.b
[^T6e@GfRcfb)G&M]XBT3@6_CeX8f3_B<M;gT<,\^cW72)7:>MBTa^I8/Aeb<>:^
_A?]UVN6LEWU55fV<KD_Pd,bK.0b^&WV/4eKeH20F3HYaKe7ET0^b,?-KD8VDE/1
^d2A;4\&d^=.ZJ/+?\+1OQJaT;;[_3I4Y:I)C[DP?V[5V?Y_U@f<gT)J9WEI3;I#
D96R&dS87GL=/[[;dd>(+[G9cPJ[9L5d6=&31R9#BM_4;/W<>AC.=87@69(+8#.M
Vc=<-]TK#JAOc/(=<0XF7a&bV3J@d^Z(gBJFHgS>Oe3V&I0GBZgJ3B[e_/@XF+WF
[KF,A?Y+5OL?,_0AISMZ]IC0]7M[),?V.UUWNF(bgT@FZcdWL?(X9@?4/D=ASV<>
?b_\&ZFI8;XX[:Z4;\-H?1]IH8aS=D<J;d-Pc>gA4KA__)d)9&N)2KNHD[Qf]7Se
XgH7L]a07Ra@R]QP>R8]K81+E;8.NHI]?1B+Y-#Ea8KAMY6)c;H=PJ(bVKGe#_S5
(J2)[VC_W)-^Q@b5#;ec+-X_(DcN<]c92,8VV#-WHB0bM@J52KC>)/79ICS2&G/M
>P8T9GGBgRf0Q_]=\H#&d^)-X?B,-2PM0Bg/a^M&Nf9&[O8-Pc\[G[36/J\dC&Ed
[24=E;W/5XP9\8P;JDZ6<MULTH#:R;BE,X(Z@(>O#g6.6J5:g]8g+5I_Ze4TS6+O
0A?EA5RP/2[VZ02_V?NDV-AD0d^PH_[>/3./XT4G=(dZ:].+5+<SE_R518O8-?2^
OC\-W3H^-L:QRIc&/&f(0.DF/[g0_3<F&94#P&=Y)UF0?a&ZD\(6X9f5&b,GdR+O
Z3]\T/9H;IU=JTf+b[+K->E]7)DeZLKY-]XG<[QMK_eLPE,MfZ7INXQ1]<UIgfRN
RZ&P?cZSfWQ?N-@:GCBUSB#;R1).Mf>M7Gb?C]G&(cb8XDB+Y_9Rbc#e;/_4XY&X
J\^)G.0[1):0[PUI__Pg76[\FP4F=B7\>DBR-TZ=#COCgH-UY7J]J9dR80(dK686
b:Z\PVT_+b[0DWZ5gRKD([,eC12LXUDF>>ZfXI4IKGPBTVVf9S7YN;G+R)3>P&8#
07PUW<a:9Ua3QE6MfWTf6@dS\=.7aP>FF(L&+,F.V:+(,gOg]:Af))#8HNYIeF.9
&CH])7\HVeOdY_[FR:+_:9QgY.2Ca.]D3HI6462NPLV;@Y/+D2_T>]?W+[@.]M8f
E(A^UdHZ\deNHAQLN-J;39S^EDXGU6b(\cL[=4=9^,YJSf+S]/SQ/.8YeC2B@97P
Kc12Y&]FNT@19BHMgSV(DLW:ZVg(&LWC[ag]3B1MOK27+0#G+<HJD\?-a1#/,J1-
I;V:PFM9b0^8@G4U/YLG-[Z57(OPgS>gF9;;>PM..U-\H788H:ETU;>VB3&1A6a[
g8X[38+Y-W8AN3JQ182GWSVH=T?QbN4dUf<dO6a1UE2R&^^G4g@:R7^EWbUXYO^M
F^TSM<O<-#/(/=)\(?bF9NT/c3d4E\\Me?0<RAHfHH0:KO+4[Ub^d6-ZSf]aH,==
?,D=:X6ZdeX272U\&Q.N>0b,J&@ON?VRcQ8\ISc6)Aag6eT0[_@P;8<eF6=-AU4/
>+O#V0bMaVb4eePS,5L(Q.d[c=Q&\aPYVeM7/G4_Me4RN0;af,;/0Eb\=<#RZA+1
N&:85gLZY1YaOI?L=bH#g>PVVT,c(V+CA5OVSIS9+6\Zg#G@7I/TVH_L9Vfa0\T0
M+KZaFR3;e.V@VS;^DX4O_>N<N7<0Y13Vff1Mc26YUXL91U8+[<6AJ<(RX)Pa?4W
0V:UFP<+K28F\-c\)#;5]LeMK.TcaE_GM-BZF,E1;aZPE(A&bILe@\:L?\b_=X1_
O&370a/Q897K56R:0HgI<2[G&:R3bU>ad<HMK.0KbK<8G6P]VJ(bP)O^Ie#I,)(N
WM5Ae1b72Cd,0?.K8F^6<8aMC,DYXaA\X>a.)KO]a#L<7=W<S/f5<0+3(Yg?P.[:
WU9;P<1Z:W5\/JHSdEf51-EEBY<AFHT#<=>=8OL>bN=J>9/_SHONQ-WEC=58L\dC
83TCOW4JTGU4&22gY^e=8fXM-OGbI)JcSM,94[(3gcfGf46fYOT?LFFU^8WEEZ7.
9SQ[[SV]G<[QYEU7<H\d8U?Xc@]>f;fHBH5,=V?M5FTH)RK<_8fG=E;9Q6,aS\11
<\+P[SYH433ZJ.)O?X\7_g4d5XcQ>H0P\J5MT8<Qgd&71cMdaJ]@I;De6KP59;L6
76OELWO(547MQ<e<@[OD7RW&TW/^6/La&VP[MOUM@;2@KB-(S4<X5NT4)Xc(41VH
L<^,F]TMW<5d(:d9c/a=bG7#a)OI]1HSd3gF@e^:&@#XeN4S30d?>03VW><Ycb)&
(]MPMC6(9QS0DO,CODD::[R<L_1;MLJKLgI3W2N.1\Y5W?O01BEO:)ATL0S<7eeV
R.&QW@Hg29Kf4^2SdF1Bg6H[AEF]7?;-]\5>.#MS]b)F_QYTTgK^@Fa]6]VX.6_K
>J07E<6Ec]8FJQ,ZV7V\\1L:OC6M2ReRXO()A634c0O@F(DPOQ:G(b4_?DfWZ#;A
)fSRZYH(R[1^V83IMUfdU,B]PK@4;<c0bLfYe8O3CULe2XGd0f_=g<f&6<@GMN=6
7Ked/H6EePE;]1&DH#5aK)K9:aWK=bZ)@:@5(O?O#G9U#IXdI3U&<>>F>#;JV-(.
5K<13V8gbOYf2QWLML:AJb?L&9<V#PC/+[K1PY5dK;^f&-9Nab7E>cf:b808[V&e
E)=,WXXRWB:NA7D3S=P@;IUa7UdI6C/\ZMOQB0>(dBBU7g1^;BR)G\dOM[ce2_=d
716H&XX\Ug9L=J:N)/RN=fWE.9BR;a9U6==1#S2)&9@30c0UO;M+TGQ/=5P)_>C2
R?c4[Ld6U(R4Df^OHcAGWf.)UfJN>.DZI51(\1DJO(OKf,C/+A&5cBMZ(gI]5)aH
eaFP02L)LVEBRA&/WRA=W7dH:Oc_a1b6N)R-_IX2UE?+RRacHZ[[41N_T7J0JLNP
Z+6817X6bN,A#D>0+0D0JG)(3d55dEV9E4YQ;b(J90f\df-DDa\dK:TN&ONL/E-C
QLcYb]d=#_^0Z4be(_SP@f?->+AA><.IJ,?S<bI>)<JJE)f98))Q1Y^,-P#>4\e/
=b_-PP;d15ZPcIOaGX32G<S5P@Hb5c;F9@J_ZU0Ba?(HX[D5\19)HC>0Jbg8/C\\
@^Z&RLD@ADcBN)ed:YQ#D4/JcUbQU[ZT<88)W>4@F1:IGSPa.>>7WdQBdYD3I9HF
VBN3ZdKDO)4:X4b)O&RPA0O?T0.;S]113BUYA^d8]=.dHMLGQHUgg)T8MZ_=6WLf
c.Je(&N(^1PEAUgL61c>6F8KT1Q5_8DSfA4c8(1;.S&PR/LfMZ@8Qe4&^QEDU..X
[egN_@5WZTQfEUUFG.d\MK@SWHdGH;A9f]U86VEOH:-O3AZ<0)cZ9J=]]M0PIB=f
K=T4EI/T3)Q<d4_ERRF<HT_FNUd,-)5KRaA6LOGB?=3>,SM>H-KKEHLK@ULcdbc&
;&R(89GNAD<c5Rg[;G^KS#4]&:(UAcXT083,GQ(T-a]?<+8bEV4>6S[QMCXQWB7C
N5S#AaWTcVSZJ9I2O.b_/PB.NWK(f9]KG\#[H@P&BDX;WGcI[,XWU,=K0QOF)gUP
PUENa7.A;8?+VR;8)Q3LWdgS2gD)Q933;OE]1IY@g1,=V.N>Q5PQVRTUK<_JNDRR
AVb86cI=_WU=CT&;X;O2VU)-\J/41.a=Z@(.WM0MX&52PFOdVb5fRH:dGggV(=?S
K4?+Gb[RP^(gO-TY^fdA4H=][#[Q+7]=cP#O1gb<C3KO2<VRNU4e]U^E7GV/F7(H
0SRA\?HYHfCd_SX?;8L=K]\&AQefbF<<c8_B@@9f6(92^KM@W#3;R/gUUQRGFN/8
(CWf<F/gC^e)dN:c+e--V_JFLZ7T7Qac3W21,=^O(^2@^>)NKHXT9C]C][U9QQ>8
NG]83UXCDO@eHW00-^QCf>We)FW&72T7FP-.<gS&Q\NYdg<49H#9b3#&-;L<TBSE
FLRHY_+b>.CR&;2Qe=C35g2ZO87.?4O[G/>OT;^@&TRga5I5WO4QIGC>XD@aSa0O
70&a6#]T)N@;VGBgJEdF9S^1)ZH9\2S/MLW&9SBO3R^1.,C+b@)[P??[g^RA#)c>
#3f#&WeV?D=A\]@7^OJ04/2KbOE^?>c(&NQML,)c<A]:YB]&Y<Y-5fJ&e]TCQOe^
]Ea\\-@(K\EY:H>)\afTZ((8E,Y?\-[[aDd<9OYa4\PeT<MN@],FU:geQbKdHf.I
L8FH=NVLcE161?8QV+)cg0aX-?\1ReO3M#=\N&FZb/BBDGe//H\KH_fR4fP+5=\3
;_T5eHDcOKO]</#S-f7b:+U1B,D=cCP:[BP0V/M1^MaXWPC(4H;e7H(J[+RfNP=B
L&/VS2E&JL>2BOA4[MOSFM;D;[#<<RKA.H:HC&O\VUKS<L)-7(Lac7E:8V7fBBGU
PXK(UH7?<BbM=&<Cf=1Y];,YTE\LNQW^0ZYgg(0+3KX^UMdO^()JPJG/6>cKZR-N
5aP88CW]5;.]ZH\\cP+_7URg)+@=6VJ-TLL1RNS0VY?9K+X+a(gP[^[O@bRBR.&Y
:NF^FZSHf=V>N\SS8K>eX=P\[V?15RCZWUL)NW):O:>ORI)aX5?&aa61Q?31^FW7
g0JK3&WDRFafZE_f(Z5=-=EN[;\L3eY.XIT(E00OF=]A)H,^Pg_EQVVL(_@K?e.L
TXLS^LGJaIX57KZ6&MH1CC7eX5fKZdc1I81UUfdGCX&X&(47f(d+.5BTd[R+fG[;
.;XA)-a#G^C:O13J8UR+E4-C6VL47&#-BKVN9HC@fL5<A74YT@@BXFF_7EGO=aUI
]CMc9XRF)Ff#+<G]5@#b.SJMXZ0\PfF9ST=ZD/CC>@Y;#4U.J#DDYcd1UDTN-MKD
7&S9N,JEKeSR)OPIF2YH1c]ER=BV+8BPZ:(+Z43(>a29;4B0<R#)2Eb.^BA8W8BA
?98W1:J&)X(Z9>J^EDg&<Zb+d8SY3.@W2>&YaK@@Z3,@M6/AX@6cc[C8AEMB?S_R
[^I>HXOf/DB5;P9EW?JXRJgbQJVO7PO@&C6-R7L;G<A//D2KVVPg@FE4fU#\2LcO
eaLG_Y\B<eK@RP1]/CP:Xcf,]O03MLX#+2dVe[SPcE[3a).cY^)GI3Nd+EM+8^f3
01>MaGX2RQRUM>P;Y\P3=-7GRc7<_OY#5@K=&?M[^]=M]I>0_518U_9<7ZNEC>\5
;@Re_Kb9E3e75SMMR6BYZ,IZSJQ>34.KfOJ,dV:@DOQX0,g&S(01A5;?BgG@(c06
2;?@c<WY(PRb]EK+JF6.K@R9ITT;[O]Z)5A]=AH?W_F8:eg.,TJAf.1=aGYgHGL1
UH9_QZ/G<AdI0d4H697A\L&712dU4)A;dFaD-UM+Xc>P(AKVgS3,6I-cM1JaZ9F;
OB)5.Yg(U76A<2TV[,04;DZTZf-XG+3.)=bY3P==_RRV3H4=4TYLeL#2e0<ZOD)f
C[8Fb\9>1]X+5+9J^>:N;1FcXCa,2+SQXc+A;XRHNg)_cZ>JT+]VeXaBUIbcPR0G
?7[@;E:Dc0.D3O^+UW@e>/1Aaf5QH#PPAadXPNIQZW<_d=0_\HNE#)5R=^1HF=T-
6S<FGZ5J9G59=-<WF=e6JOc(?9#eB1QH-8,a?,8/>-(9X[Q#U11I;FgAYX)/_cNJ
-4DGV\SDY,#;2_=;N#I^K:B&^4cfcQAW+I;LDdHGRP)PQJ+(2aaLaS<RA>c9^31<
0>3]g6d?dcVUK:fXC[SZ>.I);gW;#c_c\RJ>1MV;Wd/eNA3c#d1/.^cJc+e?^0H_
2-O5/0\,Ig40f2-3^>E.aOT0,@:U^KUg^HQbbAdB&a]0+DN7Q3QS7g#]+DI\<e)6
@LZ/1V,YbJRa13Q&aX#L2#FQ7H<.G/;?I(C-YZS<.3ENN1I3_^L#(3H,cU:9<f_:
<6Rg4>.R^<_O3SZ>,HH?L3IDT7AU\B7F#5b6K0Kg3N_9\7;T@@]-P@[a^Q9ePUI(
5f,2^&@\;K&1/@gN[,eV8[TL4EA+E]QL+/X4Peb^H21e](ZgB>PCVC/QCf^g:/dS
DYX8HME=[A)^J&7\-VBM?I4/PG<81](@.Z+PfB2B]M1-N&d8LaO^J\9ecCRGE\8@
64,GcM5[ANR5^14V#?:@</J69(6Pc.=5W^[?Ig\C<>6=)K1[JFOK2d3:4V?8MXYf
aPcGN.D^f]M7ed>_Tff(KV);M.W7SD0^LD93+X(,7DY]f2(+LcTT<GKK<>1:L298
Z>&>&IaD\XNSS/4L)VQd&@Pd9B:aHfF8@=H8a26Z94B+fE&<JRI5WWaK3;U9g1JR
C)bO9g0f4)3;6GKLdXL1KW5:=dGgf=DQ.F/?((<QJ_Z5d^RC5^=374]<38;#@f]8
\[\3V70HC,8K>]eAEW[81->Oe@CY<\fW@b8[K.bf+Mc,#gMd=Z87SEW,P3K=dGe>
A3>&7TA3e8K^)5@/1)4HGR=L,6P&gTR&]b\HV?0L<GMQVH9UMTJ&cVIdN-(8+6@P
U)HSMB-1G0<;&.;IU9;bL+V>-?eJ=Zc=-_PU4X;P+]M)QEYMO5dg[,NX>BT^g1XL
f1\aB7>Z.#X]FaK<<#[:JBP@YNc/)\-:bPI@NO:cNF>aJ.gg(&>fR_Y02E=J)@gL
a.81+SPcF15I4BBXT&LRAV_4,NIKP#WV(RP,E#NAO:c_OC\<Ag01.a\]6X>KJ-f,
GV/T-I.ISd+X:+R6U]<FM]H#>P5dKG7AO^5I/XRI5:#3b9Y73ZL]LP5QU4#=>9OQ
\5#AJBCHAgK^+N,,\GVaDeG-L(W7.03Wa8S05ZbddDJY^F0MA^6M1_EUe^8R2Y#Y
B1_>F6bGP1QcIRN:Y1Qa-X@5P\-S2W5@PYdS@EF7c;RU9YR#9&=R+S1MRY0:AKTa
)\Ie2@<fPHRbR=R/^;-_2WK&O3-SOg2P2JTOZ3d+GPEg?b)8F[FVI?aWLbA\^)K&
4-YS.Og.C>JS7/65)U>c)P;Y8L#@._<.I;K\UdVdQ[2;M3=cW)fdN>@c_)7(0JXb
E8\BdG;#Aa,&?YPG@Ub]EfKFcQdMD:7LDb^fY.@gHMcY/J7U=@NR^5dDQU-M;-FO
>.7^d4[:0bKHgKa:R:^g8E/d9aQVVUCbS6<.<Y-KL?AK-E#EYgY;fX(=F6Nc4YTM
8U00N7\CXA7MY#OcQ6=54\J-CH-3A5edTgB&#K:7-(E5+/E=UEcIX2?6#1DHY<?\
V7_C9K4\;<8[J.4W8UTH]?4J>K+GPC8JPA]>B-7OD.N92S<F_[O##(A\Ie\(3/Lf
Ie^&dW<IPOV)3AS,K8ZbMNZ]I)M-04dHNd[>]D(>,eS&Z<b)^2FV[ROP\YWH.6;e
^O_-^VZ.#M8ad@EUFGH\E.OK4<.\YDVM/5+)+J&Q=8Q)3;dSS<G:DgN4X:<(,e5e
J1[N;F79F3_E9CWTUM[bKVJB6D/YDe@51.b5(3M1EN^]8;D=K9dW5_,WKPGSdL6f
SK6,SgDc7DB,4\gBT-LH2bE3g(8HSR#,&&dLBY3#_>C0>;Vb(&_g]:XM@ecI,.@L
E;T1f-7c1]DeB3[4?(S2(6#;2aG:TAX3VA(Hac1E<KQeW]4:5ZOZ]#?.LgIC/:7Y
1&N:44V>>S4&,P393^#aR+MdRVdH(+.2FOB(WI.6J5;<_(3c6YMcG2E:^]2V&\>@
DgN;NYU_#,M]FPI\;g7<)3^N)M68CVF;(G_U;7Q:[6>XR<+Y(HWQA]Qa;B6Y[JU)
B.b?B@N2+b2?S<X8fQGU:b-DYc3M_Z#/HV3TAObb9DA[L@eYH;]7P0WZ.L0JI_I0
+2F?3:J9:@9PF^&6.DS0QOOfCQa^MXCV2U_C23b2H0c-Ca3V[LYZ6>Oc)f0CM.@3
HBK0eB8[@BHT2(5[8UI&@e_1^b[H&?-6JJ][c,^C@ZZ&A(S63gH(7/G[?^]CL#E+
S:>YX8DR@(\MW56G-IYK9AP]LYHKZTN34^9D3GL=3U/+]OGUZb&fHJ+7#1;>6S41
4?D+9dFeOJM?J1ST&#6+@_\)XU@AIZRP6Je\Uc.(B8[\++^Uf(=]dg#-;/29^<:.
BJ#.;VCS6)eHC@cdf78Gd[_4<\X#Z-PL)IUBY>7R.Q;4@=3de^W10Hd>:)AI]YgV
J6MDMNMgGaR2EO#D3UW2C-3g<SCS?C26CEC.>@CR-+L4bY2;bVQ/f@&).QX;Ua5]
<OL_..N-+7Q\gZ1T6,W<5ENH/2<ET831,WI#3,A>T5=<bD?;a[f3#:YWQ\ZN@2I:
@PI[\9eAW];?Gg7(Ya(C;#OGCP=K_bDWI=&CLeAI^cXfd3W^DgR\>([Z6XO_KOI.
aE&-;4BRHcYAE#V.2-EQSJTMYB,\C,1;PB)B;9_65)H&,-,(.0PK[C;5#;5J1I#e
[aL67E>FBU<8HK45<6QQ?JPALd-?Y-?S^MP>K>M@T8+U[>>,P+4aT(H+5>0V5+&-
TVX:5g0#)BRgD?>V=WCS9M[7KR_NVNWXF09T[dP?_VCN-86BB1A=cA8:K+2\BHER
]P_[UU:\C.^,RP0S2Af(7DX[#_f>]1b<2297&B^A\-QWgL>T=J@gP=W-E>?QU&Z-
>[>GIb]_Z\ZcDSWMR2G&b2TX7O&(=(K)K:Q+0.2T\f.,X8);b=;:H0,I9gFeN>FA
E,X&ZK1OBV6?M;C1.+/]P]9(5_(4OOTdTDQf/cB2O0N51e0<2:g\[71Qc806QEd-
(PQH2&7c4+;1?<IN@_Ub94ZI-Ce&PF&e6gF1VIDW3N@;_;]\](R@<6aNUVE<HMW3
-+&X(K[B)#X@32Q(&0J;f.,aF1.T09?F?$
`endprotected
