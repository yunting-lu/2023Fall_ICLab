# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA180_512X64X1BM1
#       Words            : 512
#       Bits             : 64
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2023/10/19 20:58:19
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA180_512X64X1BM1
CLASS BLOCK ;
FOREIGN SUMA180_512X64X1BM1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1005.020 BY 294.000 ;
SYMMETRY x y r90 ;
SITE core_5040 ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1003.900 282.580 1005.020 285.820 ;
  LAYER metal3 ;
  RECT 1003.900 282.580 1005.020 285.820 ;
  LAYER metal2 ;
  RECT 1003.900 282.580 1005.020 285.820 ;
  LAYER metal1 ;
  RECT 1003.900 282.580 1005.020 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 274.740 1005.020 277.980 ;
  LAYER metal3 ;
  RECT 1003.900 274.740 1005.020 277.980 ;
  LAYER metal2 ;
  RECT 1003.900 274.740 1005.020 277.980 ;
  LAYER metal1 ;
  RECT 1003.900 274.740 1005.020 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 266.900 1005.020 270.140 ;
  LAYER metal3 ;
  RECT 1003.900 266.900 1005.020 270.140 ;
  LAYER metal2 ;
  RECT 1003.900 266.900 1005.020 270.140 ;
  LAYER metal1 ;
  RECT 1003.900 266.900 1005.020 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 259.060 1005.020 262.300 ;
  LAYER metal3 ;
  RECT 1003.900 259.060 1005.020 262.300 ;
  LAYER metal2 ;
  RECT 1003.900 259.060 1005.020 262.300 ;
  LAYER metal1 ;
  RECT 1003.900 259.060 1005.020 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 251.220 1005.020 254.460 ;
  LAYER metal3 ;
  RECT 1003.900 251.220 1005.020 254.460 ;
  LAYER metal2 ;
  RECT 1003.900 251.220 1005.020 254.460 ;
  LAYER metal1 ;
  RECT 1003.900 251.220 1005.020 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 243.380 1005.020 246.620 ;
  LAYER metal3 ;
  RECT 1003.900 243.380 1005.020 246.620 ;
  LAYER metal2 ;
  RECT 1003.900 243.380 1005.020 246.620 ;
  LAYER metal1 ;
  RECT 1003.900 243.380 1005.020 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 204.180 1005.020 207.420 ;
  LAYER metal3 ;
  RECT 1003.900 204.180 1005.020 207.420 ;
  LAYER metal2 ;
  RECT 1003.900 204.180 1005.020 207.420 ;
  LAYER metal1 ;
  RECT 1003.900 204.180 1005.020 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 196.340 1005.020 199.580 ;
  LAYER metal3 ;
  RECT 1003.900 196.340 1005.020 199.580 ;
  LAYER metal2 ;
  RECT 1003.900 196.340 1005.020 199.580 ;
  LAYER metal1 ;
  RECT 1003.900 196.340 1005.020 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 188.500 1005.020 191.740 ;
  LAYER metal3 ;
  RECT 1003.900 188.500 1005.020 191.740 ;
  LAYER metal2 ;
  RECT 1003.900 188.500 1005.020 191.740 ;
  LAYER metal1 ;
  RECT 1003.900 188.500 1005.020 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 180.660 1005.020 183.900 ;
  LAYER metal3 ;
  RECT 1003.900 180.660 1005.020 183.900 ;
  LAYER metal2 ;
  RECT 1003.900 180.660 1005.020 183.900 ;
  LAYER metal1 ;
  RECT 1003.900 180.660 1005.020 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 172.820 1005.020 176.060 ;
  LAYER metal3 ;
  RECT 1003.900 172.820 1005.020 176.060 ;
  LAYER metal2 ;
  RECT 1003.900 172.820 1005.020 176.060 ;
  LAYER metal1 ;
  RECT 1003.900 172.820 1005.020 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 164.980 1005.020 168.220 ;
  LAYER metal3 ;
  RECT 1003.900 164.980 1005.020 168.220 ;
  LAYER metal2 ;
  RECT 1003.900 164.980 1005.020 168.220 ;
  LAYER metal1 ;
  RECT 1003.900 164.980 1005.020 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 125.780 1005.020 129.020 ;
  LAYER metal3 ;
  RECT 1003.900 125.780 1005.020 129.020 ;
  LAYER metal2 ;
  RECT 1003.900 125.780 1005.020 129.020 ;
  LAYER metal1 ;
  RECT 1003.900 125.780 1005.020 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 117.940 1005.020 121.180 ;
  LAYER metal3 ;
  RECT 1003.900 117.940 1005.020 121.180 ;
  LAYER metal2 ;
  RECT 1003.900 117.940 1005.020 121.180 ;
  LAYER metal1 ;
  RECT 1003.900 117.940 1005.020 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 110.100 1005.020 113.340 ;
  LAYER metal3 ;
  RECT 1003.900 110.100 1005.020 113.340 ;
  LAYER metal2 ;
  RECT 1003.900 110.100 1005.020 113.340 ;
  LAYER metal1 ;
  RECT 1003.900 110.100 1005.020 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 102.260 1005.020 105.500 ;
  LAYER metal3 ;
  RECT 1003.900 102.260 1005.020 105.500 ;
  LAYER metal2 ;
  RECT 1003.900 102.260 1005.020 105.500 ;
  LAYER metal1 ;
  RECT 1003.900 102.260 1005.020 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 94.420 1005.020 97.660 ;
  LAYER metal3 ;
  RECT 1003.900 94.420 1005.020 97.660 ;
  LAYER metal2 ;
  RECT 1003.900 94.420 1005.020 97.660 ;
  LAYER metal1 ;
  RECT 1003.900 94.420 1005.020 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 86.580 1005.020 89.820 ;
  LAYER metal3 ;
  RECT 1003.900 86.580 1005.020 89.820 ;
  LAYER metal2 ;
  RECT 1003.900 86.580 1005.020 89.820 ;
  LAYER metal1 ;
  RECT 1003.900 86.580 1005.020 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 47.380 1005.020 50.620 ;
  LAYER metal3 ;
  RECT 1003.900 47.380 1005.020 50.620 ;
  LAYER metal2 ;
  RECT 1003.900 47.380 1005.020 50.620 ;
  LAYER metal1 ;
  RECT 1003.900 47.380 1005.020 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 39.540 1005.020 42.780 ;
  LAYER metal3 ;
  RECT 1003.900 39.540 1005.020 42.780 ;
  LAYER metal2 ;
  RECT 1003.900 39.540 1005.020 42.780 ;
  LAYER metal1 ;
  RECT 1003.900 39.540 1005.020 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 31.700 1005.020 34.940 ;
  LAYER metal3 ;
  RECT 1003.900 31.700 1005.020 34.940 ;
  LAYER metal2 ;
  RECT 1003.900 31.700 1005.020 34.940 ;
  LAYER metal1 ;
  RECT 1003.900 31.700 1005.020 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 23.860 1005.020 27.100 ;
  LAYER metal3 ;
  RECT 1003.900 23.860 1005.020 27.100 ;
  LAYER metal2 ;
  RECT 1003.900 23.860 1005.020 27.100 ;
  LAYER metal1 ;
  RECT 1003.900 23.860 1005.020 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 16.020 1005.020 19.260 ;
  LAYER metal3 ;
  RECT 1003.900 16.020 1005.020 19.260 ;
  LAYER metal2 ;
  RECT 1003.900 16.020 1005.020 19.260 ;
  LAYER metal1 ;
  RECT 1003.900 16.020 1005.020 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 8.180 1005.020 11.420 ;
  LAYER metal3 ;
  RECT 1003.900 8.180 1005.020 11.420 ;
  LAYER metal2 ;
  RECT 1003.900 8.180 1005.020 11.420 ;
  LAYER metal1 ;
  RECT 1003.900 8.180 1005.020 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 988.680 292.880 992.220 294.000 ;
  LAYER metal3 ;
  RECT 988.680 292.880 992.220 294.000 ;
  LAYER metal2 ;
  RECT 988.680 292.880 992.220 294.000 ;
  LAYER metal1 ;
  RECT 988.680 292.880 992.220 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 980.000 292.880 983.540 294.000 ;
  LAYER metal3 ;
  RECT 980.000 292.880 983.540 294.000 ;
  LAYER metal2 ;
  RECT 980.000 292.880 983.540 294.000 ;
  LAYER metal1 ;
  RECT 980.000 292.880 983.540 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 971.320 292.880 974.860 294.000 ;
  LAYER metal3 ;
  RECT 971.320 292.880 974.860 294.000 ;
  LAYER metal2 ;
  RECT 971.320 292.880 974.860 294.000 ;
  LAYER metal1 ;
  RECT 971.320 292.880 974.860 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 962.640 292.880 966.180 294.000 ;
  LAYER metal3 ;
  RECT 962.640 292.880 966.180 294.000 ;
  LAYER metal2 ;
  RECT 962.640 292.880 966.180 294.000 ;
  LAYER metal1 ;
  RECT 962.640 292.880 966.180 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 919.240 292.880 922.780 294.000 ;
  LAYER metal3 ;
  RECT 919.240 292.880 922.780 294.000 ;
  LAYER metal2 ;
  RECT 919.240 292.880 922.780 294.000 ;
  LAYER metal1 ;
  RECT 919.240 292.880 922.780 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 910.560 292.880 914.100 294.000 ;
  LAYER metal3 ;
  RECT 910.560 292.880 914.100 294.000 ;
  LAYER metal2 ;
  RECT 910.560 292.880 914.100 294.000 ;
  LAYER metal1 ;
  RECT 910.560 292.880 914.100 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 901.880 292.880 905.420 294.000 ;
  LAYER metal3 ;
  RECT 901.880 292.880 905.420 294.000 ;
  LAYER metal2 ;
  RECT 901.880 292.880 905.420 294.000 ;
  LAYER metal1 ;
  RECT 901.880 292.880 905.420 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 893.200 292.880 896.740 294.000 ;
  LAYER metal3 ;
  RECT 893.200 292.880 896.740 294.000 ;
  LAYER metal2 ;
  RECT 893.200 292.880 896.740 294.000 ;
  LAYER metal1 ;
  RECT 893.200 292.880 896.740 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 884.520 292.880 888.060 294.000 ;
  LAYER metal3 ;
  RECT 884.520 292.880 888.060 294.000 ;
  LAYER metal2 ;
  RECT 884.520 292.880 888.060 294.000 ;
  LAYER metal1 ;
  RECT 884.520 292.880 888.060 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 875.840 292.880 879.380 294.000 ;
  LAYER metal3 ;
  RECT 875.840 292.880 879.380 294.000 ;
  LAYER metal2 ;
  RECT 875.840 292.880 879.380 294.000 ;
  LAYER metal1 ;
  RECT 875.840 292.880 879.380 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 832.440 292.880 835.980 294.000 ;
  LAYER metal3 ;
  RECT 832.440 292.880 835.980 294.000 ;
  LAYER metal2 ;
  RECT 832.440 292.880 835.980 294.000 ;
  LAYER metal1 ;
  RECT 832.440 292.880 835.980 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 823.760 292.880 827.300 294.000 ;
  LAYER metal3 ;
  RECT 823.760 292.880 827.300 294.000 ;
  LAYER metal2 ;
  RECT 823.760 292.880 827.300 294.000 ;
  LAYER metal1 ;
  RECT 823.760 292.880 827.300 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 815.080 292.880 818.620 294.000 ;
  LAYER metal3 ;
  RECT 815.080 292.880 818.620 294.000 ;
  LAYER metal2 ;
  RECT 815.080 292.880 818.620 294.000 ;
  LAYER metal1 ;
  RECT 815.080 292.880 818.620 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 806.400 292.880 809.940 294.000 ;
  LAYER metal3 ;
  RECT 806.400 292.880 809.940 294.000 ;
  LAYER metal2 ;
  RECT 806.400 292.880 809.940 294.000 ;
  LAYER metal1 ;
  RECT 806.400 292.880 809.940 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 797.720 292.880 801.260 294.000 ;
  LAYER metal3 ;
  RECT 797.720 292.880 801.260 294.000 ;
  LAYER metal2 ;
  RECT 797.720 292.880 801.260 294.000 ;
  LAYER metal1 ;
  RECT 797.720 292.880 801.260 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 789.040 292.880 792.580 294.000 ;
  LAYER metal3 ;
  RECT 789.040 292.880 792.580 294.000 ;
  LAYER metal2 ;
  RECT 789.040 292.880 792.580 294.000 ;
  LAYER metal1 ;
  RECT 789.040 292.880 792.580 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 745.640 292.880 749.180 294.000 ;
  LAYER metal3 ;
  RECT 745.640 292.880 749.180 294.000 ;
  LAYER metal2 ;
  RECT 745.640 292.880 749.180 294.000 ;
  LAYER metal1 ;
  RECT 745.640 292.880 749.180 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 736.960 292.880 740.500 294.000 ;
  LAYER metal3 ;
  RECT 736.960 292.880 740.500 294.000 ;
  LAYER metal2 ;
  RECT 736.960 292.880 740.500 294.000 ;
  LAYER metal1 ;
  RECT 736.960 292.880 740.500 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 728.280 292.880 731.820 294.000 ;
  LAYER metal3 ;
  RECT 728.280 292.880 731.820 294.000 ;
  LAYER metal2 ;
  RECT 728.280 292.880 731.820 294.000 ;
  LAYER metal1 ;
  RECT 728.280 292.880 731.820 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 719.600 292.880 723.140 294.000 ;
  LAYER metal3 ;
  RECT 719.600 292.880 723.140 294.000 ;
  LAYER metal2 ;
  RECT 719.600 292.880 723.140 294.000 ;
  LAYER metal1 ;
  RECT 719.600 292.880 723.140 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 710.920 292.880 714.460 294.000 ;
  LAYER metal3 ;
  RECT 710.920 292.880 714.460 294.000 ;
  LAYER metal2 ;
  RECT 710.920 292.880 714.460 294.000 ;
  LAYER metal1 ;
  RECT 710.920 292.880 714.460 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.240 292.880 705.780 294.000 ;
  LAYER metal3 ;
  RECT 702.240 292.880 705.780 294.000 ;
  LAYER metal2 ;
  RECT 702.240 292.880 705.780 294.000 ;
  LAYER metal1 ;
  RECT 702.240 292.880 705.780 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 658.840 292.880 662.380 294.000 ;
  LAYER metal3 ;
  RECT 658.840 292.880 662.380 294.000 ;
  LAYER metal2 ;
  RECT 658.840 292.880 662.380 294.000 ;
  LAYER metal1 ;
  RECT 658.840 292.880 662.380 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 650.160 292.880 653.700 294.000 ;
  LAYER metal3 ;
  RECT 650.160 292.880 653.700 294.000 ;
  LAYER metal2 ;
  RECT 650.160 292.880 653.700 294.000 ;
  LAYER metal1 ;
  RECT 650.160 292.880 653.700 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 641.480 292.880 645.020 294.000 ;
  LAYER metal3 ;
  RECT 641.480 292.880 645.020 294.000 ;
  LAYER metal2 ;
  RECT 641.480 292.880 645.020 294.000 ;
  LAYER metal1 ;
  RECT 641.480 292.880 645.020 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 632.800 292.880 636.340 294.000 ;
  LAYER metal3 ;
  RECT 632.800 292.880 636.340 294.000 ;
  LAYER metal2 ;
  RECT 632.800 292.880 636.340 294.000 ;
  LAYER metal1 ;
  RECT 632.800 292.880 636.340 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 624.120 292.880 627.660 294.000 ;
  LAYER metal3 ;
  RECT 624.120 292.880 627.660 294.000 ;
  LAYER metal2 ;
  RECT 624.120 292.880 627.660 294.000 ;
  LAYER metal1 ;
  RECT 624.120 292.880 627.660 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 615.440 292.880 618.980 294.000 ;
  LAYER metal3 ;
  RECT 615.440 292.880 618.980 294.000 ;
  LAYER metal2 ;
  RECT 615.440 292.880 618.980 294.000 ;
  LAYER metal1 ;
  RECT 615.440 292.880 618.980 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 572.040 292.880 575.580 294.000 ;
  LAYER metal3 ;
  RECT 572.040 292.880 575.580 294.000 ;
  LAYER metal2 ;
  RECT 572.040 292.880 575.580 294.000 ;
  LAYER metal1 ;
  RECT 572.040 292.880 575.580 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 563.360 292.880 566.900 294.000 ;
  LAYER metal3 ;
  RECT 563.360 292.880 566.900 294.000 ;
  LAYER metal2 ;
  RECT 563.360 292.880 566.900 294.000 ;
  LAYER metal1 ;
  RECT 563.360 292.880 566.900 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 554.680 292.880 558.220 294.000 ;
  LAYER metal3 ;
  RECT 554.680 292.880 558.220 294.000 ;
  LAYER metal2 ;
  RECT 554.680 292.880 558.220 294.000 ;
  LAYER metal1 ;
  RECT 554.680 292.880 558.220 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.000 292.880 549.540 294.000 ;
  LAYER metal3 ;
  RECT 546.000 292.880 549.540 294.000 ;
  LAYER metal2 ;
  RECT 546.000 292.880 549.540 294.000 ;
  LAYER metal1 ;
  RECT 546.000 292.880 549.540 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 292.880 540.860 294.000 ;
  LAYER metal3 ;
  RECT 537.320 292.880 540.860 294.000 ;
  LAYER metal2 ;
  RECT 537.320 292.880 540.860 294.000 ;
  LAYER metal1 ;
  RECT 537.320 292.880 540.860 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 292.880 532.180 294.000 ;
  LAYER metal3 ;
  RECT 528.640 292.880 532.180 294.000 ;
  LAYER metal2 ;
  RECT 528.640 292.880 532.180 294.000 ;
  LAYER metal1 ;
  RECT 528.640 292.880 532.180 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 292.880 488.780 294.000 ;
  LAYER metal3 ;
  RECT 485.240 292.880 488.780 294.000 ;
  LAYER metal2 ;
  RECT 485.240 292.880 488.780 294.000 ;
  LAYER metal1 ;
  RECT 485.240 292.880 488.780 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 292.880 480.100 294.000 ;
  LAYER metal3 ;
  RECT 476.560 292.880 480.100 294.000 ;
  LAYER metal2 ;
  RECT 476.560 292.880 480.100 294.000 ;
  LAYER metal1 ;
  RECT 476.560 292.880 480.100 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 292.880 471.420 294.000 ;
  LAYER metal3 ;
  RECT 467.880 292.880 471.420 294.000 ;
  LAYER metal2 ;
  RECT 467.880 292.880 471.420 294.000 ;
  LAYER metal1 ;
  RECT 467.880 292.880 471.420 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 292.880 462.740 294.000 ;
  LAYER metal3 ;
  RECT 459.200 292.880 462.740 294.000 ;
  LAYER metal2 ;
  RECT 459.200 292.880 462.740 294.000 ;
  LAYER metal1 ;
  RECT 459.200 292.880 462.740 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 292.880 454.060 294.000 ;
  LAYER metal3 ;
  RECT 450.520 292.880 454.060 294.000 ;
  LAYER metal2 ;
  RECT 450.520 292.880 454.060 294.000 ;
  LAYER metal1 ;
  RECT 450.520 292.880 454.060 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 292.880 445.380 294.000 ;
  LAYER metal3 ;
  RECT 441.840 292.880 445.380 294.000 ;
  LAYER metal2 ;
  RECT 441.840 292.880 445.380 294.000 ;
  LAYER metal1 ;
  RECT 441.840 292.880 445.380 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 292.880 401.980 294.000 ;
  LAYER metal3 ;
  RECT 398.440 292.880 401.980 294.000 ;
  LAYER metal2 ;
  RECT 398.440 292.880 401.980 294.000 ;
  LAYER metal1 ;
  RECT 398.440 292.880 401.980 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 292.880 393.300 294.000 ;
  LAYER metal3 ;
  RECT 389.760 292.880 393.300 294.000 ;
  LAYER metal2 ;
  RECT 389.760 292.880 393.300 294.000 ;
  LAYER metal1 ;
  RECT 389.760 292.880 393.300 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 292.880 384.620 294.000 ;
  LAYER metal3 ;
  RECT 381.080 292.880 384.620 294.000 ;
  LAYER metal2 ;
  RECT 381.080 292.880 384.620 294.000 ;
  LAYER metal1 ;
  RECT 381.080 292.880 384.620 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 292.880 375.940 294.000 ;
  LAYER metal3 ;
  RECT 372.400 292.880 375.940 294.000 ;
  LAYER metal2 ;
  RECT 372.400 292.880 375.940 294.000 ;
  LAYER metal1 ;
  RECT 372.400 292.880 375.940 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 292.880 367.260 294.000 ;
  LAYER metal3 ;
  RECT 363.720 292.880 367.260 294.000 ;
  LAYER metal2 ;
  RECT 363.720 292.880 367.260 294.000 ;
  LAYER metal1 ;
  RECT 363.720 292.880 367.260 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 292.880 358.580 294.000 ;
  LAYER metal3 ;
  RECT 355.040 292.880 358.580 294.000 ;
  LAYER metal2 ;
  RECT 355.040 292.880 358.580 294.000 ;
  LAYER metal1 ;
  RECT 355.040 292.880 358.580 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER metal3 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER metal2 ;
  RECT 311.640 292.880 315.180 294.000 ;
  LAYER metal1 ;
  RECT 311.640 292.880 315.180 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER metal3 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER metal2 ;
  RECT 302.960 292.880 306.500 294.000 ;
  LAYER metal1 ;
  RECT 302.960 292.880 306.500 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER metal3 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER metal2 ;
  RECT 294.280 292.880 297.820 294.000 ;
  LAYER metal1 ;
  RECT 294.280 292.880 297.820 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER metal3 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER metal2 ;
  RECT 285.600 292.880 289.140 294.000 ;
  LAYER metal1 ;
  RECT 285.600 292.880 289.140 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER metal3 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER metal2 ;
  RECT 276.920 292.880 280.460 294.000 ;
  LAYER metal1 ;
  RECT 276.920 292.880 280.460 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER metal3 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER metal2 ;
  RECT 268.240 292.880 271.780 294.000 ;
  LAYER metal1 ;
  RECT 268.240 292.880 271.780 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER metal3 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER metal2 ;
  RECT 224.840 292.880 228.380 294.000 ;
  LAYER metal1 ;
  RECT 224.840 292.880 228.380 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER metal3 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER metal2 ;
  RECT 216.160 292.880 219.700 294.000 ;
  LAYER metal1 ;
  RECT 216.160 292.880 219.700 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER metal3 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER metal2 ;
  RECT 207.480 292.880 211.020 294.000 ;
  LAYER metal1 ;
  RECT 207.480 292.880 211.020 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER metal3 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER metal2 ;
  RECT 198.800 292.880 202.340 294.000 ;
  LAYER metal1 ;
  RECT 198.800 292.880 202.340 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER metal3 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER metal2 ;
  RECT 190.120 292.880 193.660 294.000 ;
  LAYER metal1 ;
  RECT 190.120 292.880 193.660 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER metal3 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER metal2 ;
  RECT 181.440 292.880 184.980 294.000 ;
  LAYER metal1 ;
  RECT 181.440 292.880 184.980 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER metal3 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER metal2 ;
  RECT 138.040 292.880 141.580 294.000 ;
  LAYER metal1 ;
  RECT 138.040 292.880 141.580 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER metal3 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER metal2 ;
  RECT 129.360 292.880 132.900 294.000 ;
  LAYER metal1 ;
  RECT 129.360 292.880 132.900 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER metal3 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER metal2 ;
  RECT 120.680 292.880 124.220 294.000 ;
  LAYER metal1 ;
  RECT 120.680 292.880 124.220 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER metal3 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER metal2 ;
  RECT 112.000 292.880 115.540 294.000 ;
  LAYER metal1 ;
  RECT 112.000 292.880 115.540 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER metal3 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER metal2 ;
  RECT 103.320 292.880 106.860 294.000 ;
  LAYER metal1 ;
  RECT 103.320 292.880 106.860 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER metal3 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER metal2 ;
  RECT 94.640 292.880 98.180 294.000 ;
  LAYER metal1 ;
  RECT 94.640 292.880 98.180 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER metal3 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER metal2 ;
  RECT 51.240 292.880 54.780 294.000 ;
  LAYER metal1 ;
  RECT 51.240 292.880 54.780 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER metal3 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER metal2 ;
  RECT 42.560 292.880 46.100 294.000 ;
  LAYER metal1 ;
  RECT 42.560 292.880 46.100 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER metal3 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER metal2 ;
  RECT 33.880 292.880 37.420 294.000 ;
  LAYER metal1 ;
  RECT 33.880 292.880 37.420 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER metal3 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER metal2 ;
  RECT 25.200 292.880 28.740 294.000 ;
  LAYER metal1 ;
  RECT 25.200 292.880 28.740 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER metal3 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER metal2 ;
  RECT 16.520 292.880 20.060 294.000 ;
  LAYER metal1 ;
  RECT 16.520 292.880 20.060 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER metal3 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER metal2 ;
  RECT 7.840 292.880 11.380 294.000 ;
  LAYER metal1 ;
  RECT 7.840 292.880 11.380 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 985.580 0.000 989.120 1.120 ;
  LAYER metal3 ;
  RECT 985.580 0.000 989.120 1.120 ;
  LAYER metal2 ;
  RECT 985.580 0.000 989.120 1.120 ;
  LAYER metal1 ;
  RECT 985.580 0.000 989.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 963.880 0.000 967.420 1.120 ;
  LAYER metal3 ;
  RECT 963.880 0.000 967.420 1.120 ;
  LAYER metal2 ;
  RECT 963.880 0.000 967.420 1.120 ;
  LAYER metal1 ;
  RECT 963.880 0.000 967.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 942.180 0.000 945.720 1.120 ;
  LAYER metal3 ;
  RECT 942.180 0.000 945.720 1.120 ;
  LAYER metal2 ;
  RECT 942.180 0.000 945.720 1.120 ;
  LAYER metal1 ;
  RECT 942.180 0.000 945.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 915.520 0.000 919.060 1.120 ;
  LAYER metal3 ;
  RECT 915.520 0.000 919.060 1.120 ;
  LAYER metal2 ;
  RECT 915.520 0.000 919.060 1.120 ;
  LAYER metal1 ;
  RECT 915.520 0.000 919.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 898.780 0.000 902.320 1.120 ;
  LAYER metal3 ;
  RECT 898.780 0.000 902.320 1.120 ;
  LAYER metal2 ;
  RECT 898.780 0.000 902.320 1.120 ;
  LAYER metal1 ;
  RECT 898.780 0.000 902.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 785.940 0.000 789.480 1.120 ;
  LAYER metal3 ;
  RECT 785.940 0.000 789.480 1.120 ;
  LAYER metal2 ;
  RECT 785.940 0.000 789.480 1.120 ;
  LAYER metal1 ;
  RECT 785.940 0.000 789.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 759.280 0.000 762.820 1.120 ;
  LAYER metal3 ;
  RECT 759.280 0.000 762.820 1.120 ;
  LAYER metal2 ;
  RECT 759.280 0.000 762.820 1.120 ;
  LAYER metal1 ;
  RECT 759.280 0.000 762.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 737.580 0.000 741.120 1.120 ;
  LAYER metal3 ;
  RECT 737.580 0.000 741.120 1.120 ;
  LAYER metal2 ;
  RECT 737.580 0.000 741.120 1.120 ;
  LAYER metal1 ;
  RECT 737.580 0.000 741.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 715.880 0.000 719.420 1.120 ;
  LAYER metal3 ;
  RECT 715.880 0.000 719.420 1.120 ;
  LAYER metal2 ;
  RECT 715.880 0.000 719.420 1.120 ;
  LAYER metal1 ;
  RECT 715.880 0.000 719.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal3 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal2 ;
  RECT 689.220 0.000 692.760 1.120 ;
  LAYER metal1 ;
  RECT 689.220 0.000 692.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 673.100 0.000 676.640 1.120 ;
  LAYER metal3 ;
  RECT 673.100 0.000 676.640 1.120 ;
  LAYER metal2 ;
  RECT 673.100 0.000 676.640 1.120 ;
  LAYER metal1 ;
  RECT 673.100 0.000 676.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.640 0.000 563.180 1.120 ;
  LAYER metal3 ;
  RECT 559.640 0.000 563.180 1.120 ;
  LAYER metal2 ;
  RECT 559.640 0.000 563.180 1.120 ;
  LAYER metal1 ;
  RECT 559.640 0.000 563.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 523.680 0.000 527.220 1.120 ;
  LAYER metal3 ;
  RECT 523.680 0.000 527.220 1.120 ;
  LAYER metal2 ;
  RECT 523.680 0.000 527.220 1.120 ;
  LAYER metal1 ;
  RECT 523.680 0.000 527.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 515.000 0.000 518.540 1.120 ;
  LAYER metal3 ;
  RECT 515.000 0.000 518.540 1.120 ;
  LAYER metal2 ;
  RECT 515.000 0.000 518.540 1.120 ;
  LAYER metal1 ;
  RECT 515.000 0.000 518.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal3 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal2 ;
  RECT 493.300 0.000 496.840 1.120 ;
  LAYER metal1 ;
  RECT 493.300 0.000 496.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER metal3 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER metal2 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER metal1 ;
  RECT 472.220 0.000 475.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 461.060 0.000 464.600 1.120 ;
  LAYER metal3 ;
  RECT 461.060 0.000 464.600 1.120 ;
  LAYER metal2 ;
  RECT 461.060 0.000 464.600 1.120 ;
  LAYER metal1 ;
  RECT 461.060 0.000 464.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal3 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal2 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal1 ;
  RECT 353.180 0.000 356.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal3 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal2 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal1 ;
  RECT 326.520 0.000 330.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER metal3 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER metal2 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER metal1 ;
  RECT 309.780 0.000 313.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1003.900 278.660 1005.020 281.900 ;
  LAYER metal3 ;
  RECT 1003.900 278.660 1005.020 281.900 ;
  LAYER metal2 ;
  RECT 1003.900 278.660 1005.020 281.900 ;
  LAYER metal1 ;
  RECT 1003.900 278.660 1005.020 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 270.820 1005.020 274.060 ;
  LAYER metal3 ;
  RECT 1003.900 270.820 1005.020 274.060 ;
  LAYER metal2 ;
  RECT 1003.900 270.820 1005.020 274.060 ;
  LAYER metal1 ;
  RECT 1003.900 270.820 1005.020 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 262.980 1005.020 266.220 ;
  LAYER metal3 ;
  RECT 1003.900 262.980 1005.020 266.220 ;
  LAYER metal2 ;
  RECT 1003.900 262.980 1005.020 266.220 ;
  LAYER metal1 ;
  RECT 1003.900 262.980 1005.020 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 255.140 1005.020 258.380 ;
  LAYER metal3 ;
  RECT 1003.900 255.140 1005.020 258.380 ;
  LAYER metal2 ;
  RECT 1003.900 255.140 1005.020 258.380 ;
  LAYER metal1 ;
  RECT 1003.900 255.140 1005.020 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 247.300 1005.020 250.540 ;
  LAYER metal3 ;
  RECT 1003.900 247.300 1005.020 250.540 ;
  LAYER metal2 ;
  RECT 1003.900 247.300 1005.020 250.540 ;
  LAYER metal1 ;
  RECT 1003.900 247.300 1005.020 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 208.100 1005.020 211.340 ;
  LAYER metal3 ;
  RECT 1003.900 208.100 1005.020 211.340 ;
  LAYER metal2 ;
  RECT 1003.900 208.100 1005.020 211.340 ;
  LAYER metal1 ;
  RECT 1003.900 208.100 1005.020 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 200.260 1005.020 203.500 ;
  LAYER metal3 ;
  RECT 1003.900 200.260 1005.020 203.500 ;
  LAYER metal2 ;
  RECT 1003.900 200.260 1005.020 203.500 ;
  LAYER metal1 ;
  RECT 1003.900 200.260 1005.020 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 192.420 1005.020 195.660 ;
  LAYER metal3 ;
  RECT 1003.900 192.420 1005.020 195.660 ;
  LAYER metal2 ;
  RECT 1003.900 192.420 1005.020 195.660 ;
  LAYER metal1 ;
  RECT 1003.900 192.420 1005.020 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 184.580 1005.020 187.820 ;
  LAYER metal3 ;
  RECT 1003.900 184.580 1005.020 187.820 ;
  LAYER metal2 ;
  RECT 1003.900 184.580 1005.020 187.820 ;
  LAYER metal1 ;
  RECT 1003.900 184.580 1005.020 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 176.740 1005.020 179.980 ;
  LAYER metal3 ;
  RECT 1003.900 176.740 1005.020 179.980 ;
  LAYER metal2 ;
  RECT 1003.900 176.740 1005.020 179.980 ;
  LAYER metal1 ;
  RECT 1003.900 176.740 1005.020 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 168.900 1005.020 172.140 ;
  LAYER metal3 ;
  RECT 1003.900 168.900 1005.020 172.140 ;
  LAYER metal2 ;
  RECT 1003.900 168.900 1005.020 172.140 ;
  LAYER metal1 ;
  RECT 1003.900 168.900 1005.020 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 129.700 1005.020 132.940 ;
  LAYER metal3 ;
  RECT 1003.900 129.700 1005.020 132.940 ;
  LAYER metal2 ;
  RECT 1003.900 129.700 1005.020 132.940 ;
  LAYER metal1 ;
  RECT 1003.900 129.700 1005.020 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 121.860 1005.020 125.100 ;
  LAYER metal3 ;
  RECT 1003.900 121.860 1005.020 125.100 ;
  LAYER metal2 ;
  RECT 1003.900 121.860 1005.020 125.100 ;
  LAYER metal1 ;
  RECT 1003.900 121.860 1005.020 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 114.020 1005.020 117.260 ;
  LAYER metal3 ;
  RECT 1003.900 114.020 1005.020 117.260 ;
  LAYER metal2 ;
  RECT 1003.900 114.020 1005.020 117.260 ;
  LAYER metal1 ;
  RECT 1003.900 114.020 1005.020 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 106.180 1005.020 109.420 ;
  LAYER metal3 ;
  RECT 1003.900 106.180 1005.020 109.420 ;
  LAYER metal2 ;
  RECT 1003.900 106.180 1005.020 109.420 ;
  LAYER metal1 ;
  RECT 1003.900 106.180 1005.020 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 98.340 1005.020 101.580 ;
  LAYER metal3 ;
  RECT 1003.900 98.340 1005.020 101.580 ;
  LAYER metal2 ;
  RECT 1003.900 98.340 1005.020 101.580 ;
  LAYER metal1 ;
  RECT 1003.900 98.340 1005.020 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 90.500 1005.020 93.740 ;
  LAYER metal3 ;
  RECT 1003.900 90.500 1005.020 93.740 ;
  LAYER metal2 ;
  RECT 1003.900 90.500 1005.020 93.740 ;
  LAYER metal1 ;
  RECT 1003.900 90.500 1005.020 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 51.300 1005.020 54.540 ;
  LAYER metal3 ;
  RECT 1003.900 51.300 1005.020 54.540 ;
  LAYER metal2 ;
  RECT 1003.900 51.300 1005.020 54.540 ;
  LAYER metal1 ;
  RECT 1003.900 51.300 1005.020 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 43.460 1005.020 46.700 ;
  LAYER metal3 ;
  RECT 1003.900 43.460 1005.020 46.700 ;
  LAYER metal2 ;
  RECT 1003.900 43.460 1005.020 46.700 ;
  LAYER metal1 ;
  RECT 1003.900 43.460 1005.020 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 35.620 1005.020 38.860 ;
  LAYER metal3 ;
  RECT 1003.900 35.620 1005.020 38.860 ;
  LAYER metal2 ;
  RECT 1003.900 35.620 1005.020 38.860 ;
  LAYER metal1 ;
  RECT 1003.900 35.620 1005.020 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 27.780 1005.020 31.020 ;
  LAYER metal3 ;
  RECT 1003.900 27.780 1005.020 31.020 ;
  LAYER metal2 ;
  RECT 1003.900 27.780 1005.020 31.020 ;
  LAYER metal1 ;
  RECT 1003.900 27.780 1005.020 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 19.940 1005.020 23.180 ;
  LAYER metal3 ;
  RECT 1003.900 19.940 1005.020 23.180 ;
  LAYER metal2 ;
  RECT 1003.900 19.940 1005.020 23.180 ;
  LAYER metal1 ;
  RECT 1003.900 19.940 1005.020 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1003.900 12.100 1005.020 15.340 ;
  LAYER metal3 ;
  RECT 1003.900 12.100 1005.020 15.340 ;
  LAYER metal2 ;
  RECT 1003.900 12.100 1005.020 15.340 ;
  LAYER metal1 ;
  RECT 1003.900 12.100 1005.020 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 993.020 292.880 996.560 294.000 ;
  LAYER metal3 ;
  RECT 993.020 292.880 996.560 294.000 ;
  LAYER metal2 ;
  RECT 993.020 292.880 996.560 294.000 ;
  LAYER metal1 ;
  RECT 993.020 292.880 996.560 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 984.340 292.880 987.880 294.000 ;
  LAYER metal3 ;
  RECT 984.340 292.880 987.880 294.000 ;
  LAYER metal2 ;
  RECT 984.340 292.880 987.880 294.000 ;
  LAYER metal1 ;
  RECT 984.340 292.880 987.880 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 975.660 292.880 979.200 294.000 ;
  LAYER metal3 ;
  RECT 975.660 292.880 979.200 294.000 ;
  LAYER metal2 ;
  RECT 975.660 292.880 979.200 294.000 ;
  LAYER metal1 ;
  RECT 975.660 292.880 979.200 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 966.980 292.880 970.520 294.000 ;
  LAYER metal3 ;
  RECT 966.980 292.880 970.520 294.000 ;
  LAYER metal2 ;
  RECT 966.980 292.880 970.520 294.000 ;
  LAYER metal1 ;
  RECT 966.980 292.880 970.520 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 923.580 292.880 927.120 294.000 ;
  LAYER metal3 ;
  RECT 923.580 292.880 927.120 294.000 ;
  LAYER metal2 ;
  RECT 923.580 292.880 927.120 294.000 ;
  LAYER metal1 ;
  RECT 923.580 292.880 927.120 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 914.900 292.880 918.440 294.000 ;
  LAYER metal3 ;
  RECT 914.900 292.880 918.440 294.000 ;
  LAYER metal2 ;
  RECT 914.900 292.880 918.440 294.000 ;
  LAYER metal1 ;
  RECT 914.900 292.880 918.440 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 906.220 292.880 909.760 294.000 ;
  LAYER metal3 ;
  RECT 906.220 292.880 909.760 294.000 ;
  LAYER metal2 ;
  RECT 906.220 292.880 909.760 294.000 ;
  LAYER metal1 ;
  RECT 906.220 292.880 909.760 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 897.540 292.880 901.080 294.000 ;
  LAYER metal3 ;
  RECT 897.540 292.880 901.080 294.000 ;
  LAYER metal2 ;
  RECT 897.540 292.880 901.080 294.000 ;
  LAYER metal1 ;
  RECT 897.540 292.880 901.080 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 888.860 292.880 892.400 294.000 ;
  LAYER metal3 ;
  RECT 888.860 292.880 892.400 294.000 ;
  LAYER metal2 ;
  RECT 888.860 292.880 892.400 294.000 ;
  LAYER metal1 ;
  RECT 888.860 292.880 892.400 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 880.180 292.880 883.720 294.000 ;
  LAYER metal3 ;
  RECT 880.180 292.880 883.720 294.000 ;
  LAYER metal2 ;
  RECT 880.180 292.880 883.720 294.000 ;
  LAYER metal1 ;
  RECT 880.180 292.880 883.720 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 836.780 292.880 840.320 294.000 ;
  LAYER metal3 ;
  RECT 836.780 292.880 840.320 294.000 ;
  LAYER metal2 ;
  RECT 836.780 292.880 840.320 294.000 ;
  LAYER metal1 ;
  RECT 836.780 292.880 840.320 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 828.100 292.880 831.640 294.000 ;
  LAYER metal3 ;
  RECT 828.100 292.880 831.640 294.000 ;
  LAYER metal2 ;
  RECT 828.100 292.880 831.640 294.000 ;
  LAYER metal1 ;
  RECT 828.100 292.880 831.640 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 819.420 292.880 822.960 294.000 ;
  LAYER metal3 ;
  RECT 819.420 292.880 822.960 294.000 ;
  LAYER metal2 ;
  RECT 819.420 292.880 822.960 294.000 ;
  LAYER metal1 ;
  RECT 819.420 292.880 822.960 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 810.740 292.880 814.280 294.000 ;
  LAYER metal3 ;
  RECT 810.740 292.880 814.280 294.000 ;
  LAYER metal2 ;
  RECT 810.740 292.880 814.280 294.000 ;
  LAYER metal1 ;
  RECT 810.740 292.880 814.280 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 802.060 292.880 805.600 294.000 ;
  LAYER metal3 ;
  RECT 802.060 292.880 805.600 294.000 ;
  LAYER metal2 ;
  RECT 802.060 292.880 805.600 294.000 ;
  LAYER metal1 ;
  RECT 802.060 292.880 805.600 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 793.380 292.880 796.920 294.000 ;
  LAYER metal3 ;
  RECT 793.380 292.880 796.920 294.000 ;
  LAYER metal2 ;
  RECT 793.380 292.880 796.920 294.000 ;
  LAYER metal1 ;
  RECT 793.380 292.880 796.920 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.980 292.880 753.520 294.000 ;
  LAYER metal3 ;
  RECT 749.980 292.880 753.520 294.000 ;
  LAYER metal2 ;
  RECT 749.980 292.880 753.520 294.000 ;
  LAYER metal1 ;
  RECT 749.980 292.880 753.520 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 741.300 292.880 744.840 294.000 ;
  LAYER metal3 ;
  RECT 741.300 292.880 744.840 294.000 ;
  LAYER metal2 ;
  RECT 741.300 292.880 744.840 294.000 ;
  LAYER metal1 ;
  RECT 741.300 292.880 744.840 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 732.620 292.880 736.160 294.000 ;
  LAYER metal3 ;
  RECT 732.620 292.880 736.160 294.000 ;
  LAYER metal2 ;
  RECT 732.620 292.880 736.160 294.000 ;
  LAYER metal1 ;
  RECT 732.620 292.880 736.160 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 723.940 292.880 727.480 294.000 ;
  LAYER metal3 ;
  RECT 723.940 292.880 727.480 294.000 ;
  LAYER metal2 ;
  RECT 723.940 292.880 727.480 294.000 ;
  LAYER metal1 ;
  RECT 723.940 292.880 727.480 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 715.260 292.880 718.800 294.000 ;
  LAYER metal3 ;
  RECT 715.260 292.880 718.800 294.000 ;
  LAYER metal2 ;
  RECT 715.260 292.880 718.800 294.000 ;
  LAYER metal1 ;
  RECT 715.260 292.880 718.800 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 706.580 292.880 710.120 294.000 ;
  LAYER metal3 ;
  RECT 706.580 292.880 710.120 294.000 ;
  LAYER metal2 ;
  RECT 706.580 292.880 710.120 294.000 ;
  LAYER metal1 ;
  RECT 706.580 292.880 710.120 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 663.180 292.880 666.720 294.000 ;
  LAYER metal3 ;
  RECT 663.180 292.880 666.720 294.000 ;
  LAYER metal2 ;
  RECT 663.180 292.880 666.720 294.000 ;
  LAYER metal1 ;
  RECT 663.180 292.880 666.720 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 654.500 292.880 658.040 294.000 ;
  LAYER metal3 ;
  RECT 654.500 292.880 658.040 294.000 ;
  LAYER metal2 ;
  RECT 654.500 292.880 658.040 294.000 ;
  LAYER metal1 ;
  RECT 654.500 292.880 658.040 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 645.820 292.880 649.360 294.000 ;
  LAYER metal3 ;
  RECT 645.820 292.880 649.360 294.000 ;
  LAYER metal2 ;
  RECT 645.820 292.880 649.360 294.000 ;
  LAYER metal1 ;
  RECT 645.820 292.880 649.360 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 637.140 292.880 640.680 294.000 ;
  LAYER metal3 ;
  RECT 637.140 292.880 640.680 294.000 ;
  LAYER metal2 ;
  RECT 637.140 292.880 640.680 294.000 ;
  LAYER metal1 ;
  RECT 637.140 292.880 640.680 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 628.460 292.880 632.000 294.000 ;
  LAYER metal3 ;
  RECT 628.460 292.880 632.000 294.000 ;
  LAYER metal2 ;
  RECT 628.460 292.880 632.000 294.000 ;
  LAYER metal1 ;
  RECT 628.460 292.880 632.000 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 619.780 292.880 623.320 294.000 ;
  LAYER metal3 ;
  RECT 619.780 292.880 623.320 294.000 ;
  LAYER metal2 ;
  RECT 619.780 292.880 623.320 294.000 ;
  LAYER metal1 ;
  RECT 619.780 292.880 623.320 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 576.380 292.880 579.920 294.000 ;
  LAYER metal3 ;
  RECT 576.380 292.880 579.920 294.000 ;
  LAYER metal2 ;
  RECT 576.380 292.880 579.920 294.000 ;
  LAYER metal1 ;
  RECT 576.380 292.880 579.920 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 567.700 292.880 571.240 294.000 ;
  LAYER metal3 ;
  RECT 567.700 292.880 571.240 294.000 ;
  LAYER metal2 ;
  RECT 567.700 292.880 571.240 294.000 ;
  LAYER metal1 ;
  RECT 567.700 292.880 571.240 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.020 292.880 562.560 294.000 ;
  LAYER metal3 ;
  RECT 559.020 292.880 562.560 294.000 ;
  LAYER metal2 ;
  RECT 559.020 292.880 562.560 294.000 ;
  LAYER metal1 ;
  RECT 559.020 292.880 562.560 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 550.340 292.880 553.880 294.000 ;
  LAYER metal3 ;
  RECT 550.340 292.880 553.880 294.000 ;
  LAYER metal2 ;
  RECT 550.340 292.880 553.880 294.000 ;
  LAYER metal1 ;
  RECT 550.340 292.880 553.880 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 292.880 545.200 294.000 ;
  LAYER metal3 ;
  RECT 541.660 292.880 545.200 294.000 ;
  LAYER metal2 ;
  RECT 541.660 292.880 545.200 294.000 ;
  LAYER metal1 ;
  RECT 541.660 292.880 545.200 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 292.880 536.520 294.000 ;
  LAYER metal3 ;
  RECT 532.980 292.880 536.520 294.000 ;
  LAYER metal2 ;
  RECT 532.980 292.880 536.520 294.000 ;
  LAYER metal1 ;
  RECT 532.980 292.880 536.520 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 292.880 493.120 294.000 ;
  LAYER metal3 ;
  RECT 489.580 292.880 493.120 294.000 ;
  LAYER metal2 ;
  RECT 489.580 292.880 493.120 294.000 ;
  LAYER metal1 ;
  RECT 489.580 292.880 493.120 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 292.880 484.440 294.000 ;
  LAYER metal3 ;
  RECT 480.900 292.880 484.440 294.000 ;
  LAYER metal2 ;
  RECT 480.900 292.880 484.440 294.000 ;
  LAYER metal1 ;
  RECT 480.900 292.880 484.440 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 292.880 475.760 294.000 ;
  LAYER metal3 ;
  RECT 472.220 292.880 475.760 294.000 ;
  LAYER metal2 ;
  RECT 472.220 292.880 475.760 294.000 ;
  LAYER metal1 ;
  RECT 472.220 292.880 475.760 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 292.880 467.080 294.000 ;
  LAYER metal3 ;
  RECT 463.540 292.880 467.080 294.000 ;
  LAYER metal2 ;
  RECT 463.540 292.880 467.080 294.000 ;
  LAYER metal1 ;
  RECT 463.540 292.880 467.080 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 292.880 458.400 294.000 ;
  LAYER metal3 ;
  RECT 454.860 292.880 458.400 294.000 ;
  LAYER metal2 ;
  RECT 454.860 292.880 458.400 294.000 ;
  LAYER metal1 ;
  RECT 454.860 292.880 458.400 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 292.880 449.720 294.000 ;
  LAYER metal3 ;
  RECT 446.180 292.880 449.720 294.000 ;
  LAYER metal2 ;
  RECT 446.180 292.880 449.720 294.000 ;
  LAYER metal1 ;
  RECT 446.180 292.880 449.720 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 292.880 406.320 294.000 ;
  LAYER metal3 ;
  RECT 402.780 292.880 406.320 294.000 ;
  LAYER metal2 ;
  RECT 402.780 292.880 406.320 294.000 ;
  LAYER metal1 ;
  RECT 402.780 292.880 406.320 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 292.880 397.640 294.000 ;
  LAYER metal3 ;
  RECT 394.100 292.880 397.640 294.000 ;
  LAYER metal2 ;
  RECT 394.100 292.880 397.640 294.000 ;
  LAYER metal1 ;
  RECT 394.100 292.880 397.640 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 292.880 388.960 294.000 ;
  LAYER metal3 ;
  RECT 385.420 292.880 388.960 294.000 ;
  LAYER metal2 ;
  RECT 385.420 292.880 388.960 294.000 ;
  LAYER metal1 ;
  RECT 385.420 292.880 388.960 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 292.880 380.280 294.000 ;
  LAYER metal3 ;
  RECT 376.740 292.880 380.280 294.000 ;
  LAYER metal2 ;
  RECT 376.740 292.880 380.280 294.000 ;
  LAYER metal1 ;
  RECT 376.740 292.880 380.280 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 292.880 371.600 294.000 ;
  LAYER metal3 ;
  RECT 368.060 292.880 371.600 294.000 ;
  LAYER metal2 ;
  RECT 368.060 292.880 371.600 294.000 ;
  LAYER metal1 ;
  RECT 368.060 292.880 371.600 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 292.880 362.920 294.000 ;
  LAYER metal3 ;
  RECT 359.380 292.880 362.920 294.000 ;
  LAYER metal2 ;
  RECT 359.380 292.880 362.920 294.000 ;
  LAYER metal1 ;
  RECT 359.380 292.880 362.920 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 292.880 319.520 294.000 ;
  LAYER metal3 ;
  RECT 315.980 292.880 319.520 294.000 ;
  LAYER metal2 ;
  RECT 315.980 292.880 319.520 294.000 ;
  LAYER metal1 ;
  RECT 315.980 292.880 319.520 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER metal3 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER metal2 ;
  RECT 307.300 292.880 310.840 294.000 ;
  LAYER metal1 ;
  RECT 307.300 292.880 310.840 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER metal3 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER metal2 ;
  RECT 298.620 292.880 302.160 294.000 ;
  LAYER metal1 ;
  RECT 298.620 292.880 302.160 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER metal3 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER metal2 ;
  RECT 289.940 292.880 293.480 294.000 ;
  LAYER metal1 ;
  RECT 289.940 292.880 293.480 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER metal3 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER metal2 ;
  RECT 281.260 292.880 284.800 294.000 ;
  LAYER metal1 ;
  RECT 281.260 292.880 284.800 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER metal3 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER metal2 ;
  RECT 272.580 292.880 276.120 294.000 ;
  LAYER metal1 ;
  RECT 272.580 292.880 276.120 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER metal3 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER metal2 ;
  RECT 229.180 292.880 232.720 294.000 ;
  LAYER metal1 ;
  RECT 229.180 292.880 232.720 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER metal3 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER metal2 ;
  RECT 220.500 292.880 224.040 294.000 ;
  LAYER metal1 ;
  RECT 220.500 292.880 224.040 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER metal3 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER metal2 ;
  RECT 211.820 292.880 215.360 294.000 ;
  LAYER metal1 ;
  RECT 211.820 292.880 215.360 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER metal3 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER metal2 ;
  RECT 203.140 292.880 206.680 294.000 ;
  LAYER metal1 ;
  RECT 203.140 292.880 206.680 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER metal3 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER metal2 ;
  RECT 194.460 292.880 198.000 294.000 ;
  LAYER metal1 ;
  RECT 194.460 292.880 198.000 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER metal3 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER metal2 ;
  RECT 185.780 292.880 189.320 294.000 ;
  LAYER metal1 ;
  RECT 185.780 292.880 189.320 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER metal3 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER metal2 ;
  RECT 142.380 292.880 145.920 294.000 ;
  LAYER metal1 ;
  RECT 142.380 292.880 145.920 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER metal3 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER metal2 ;
  RECT 133.700 292.880 137.240 294.000 ;
  LAYER metal1 ;
  RECT 133.700 292.880 137.240 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER metal3 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER metal2 ;
  RECT 125.020 292.880 128.560 294.000 ;
  LAYER metal1 ;
  RECT 125.020 292.880 128.560 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER metal3 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER metal2 ;
  RECT 116.340 292.880 119.880 294.000 ;
  LAYER metal1 ;
  RECT 116.340 292.880 119.880 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER metal3 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER metal2 ;
  RECT 107.660 292.880 111.200 294.000 ;
  LAYER metal1 ;
  RECT 107.660 292.880 111.200 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER metal3 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER metal2 ;
  RECT 98.980 292.880 102.520 294.000 ;
  LAYER metal1 ;
  RECT 98.980 292.880 102.520 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER metal3 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER metal2 ;
  RECT 55.580 292.880 59.120 294.000 ;
  LAYER metal1 ;
  RECT 55.580 292.880 59.120 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER metal3 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER metal2 ;
  RECT 46.900 292.880 50.440 294.000 ;
  LAYER metal1 ;
  RECT 46.900 292.880 50.440 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER metal3 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER metal2 ;
  RECT 38.220 292.880 41.760 294.000 ;
  LAYER metal1 ;
  RECT 38.220 292.880 41.760 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER metal3 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER metal2 ;
  RECT 29.540 292.880 33.080 294.000 ;
  LAYER metal1 ;
  RECT 29.540 292.880 33.080 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER metal3 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER metal2 ;
  RECT 20.860 292.880 24.400 294.000 ;
  LAYER metal1 ;
  RECT 20.860 292.880 24.400 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER metal3 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER metal2 ;
  RECT 12.180 292.880 15.720 294.000 ;
  LAYER metal1 ;
  RECT 12.180 292.880 15.720 294.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 993.640 0.000 997.180 1.120 ;
  LAYER metal3 ;
  RECT 993.640 0.000 997.180 1.120 ;
  LAYER metal2 ;
  RECT 993.640 0.000 997.180 1.120 ;
  LAYER metal1 ;
  RECT 993.640 0.000 997.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 971.940 0.000 975.480 1.120 ;
  LAYER metal3 ;
  RECT 971.940 0.000 975.480 1.120 ;
  LAYER metal2 ;
  RECT 971.940 0.000 975.480 1.120 ;
  LAYER metal1 ;
  RECT 971.940 0.000 975.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 955.200 0.000 958.740 1.120 ;
  LAYER metal3 ;
  RECT 955.200 0.000 958.740 1.120 ;
  LAYER metal2 ;
  RECT 955.200 0.000 958.740 1.120 ;
  LAYER metal1 ;
  RECT 955.200 0.000 958.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 928.540 0.000 932.080 1.120 ;
  LAYER metal3 ;
  RECT 928.540 0.000 932.080 1.120 ;
  LAYER metal2 ;
  RECT 928.540 0.000 932.080 1.120 ;
  LAYER metal1 ;
  RECT 928.540 0.000 932.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 907.460 0.000 911.000 1.120 ;
  LAYER metal3 ;
  RECT 907.460 0.000 911.000 1.120 ;
  LAYER metal2 ;
  RECT 907.460 0.000 911.000 1.120 ;
  LAYER metal1 ;
  RECT 907.460 0.000 911.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 794.000 0.000 797.540 1.120 ;
  LAYER metal3 ;
  RECT 794.000 0.000 797.540 1.120 ;
  LAYER metal2 ;
  RECT 794.000 0.000 797.540 1.120 ;
  LAYER metal1 ;
  RECT 794.000 0.000 797.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 772.300 0.000 775.840 1.120 ;
  LAYER metal3 ;
  RECT 772.300 0.000 775.840 1.120 ;
  LAYER metal2 ;
  RECT 772.300 0.000 775.840 1.120 ;
  LAYER metal1 ;
  RECT 772.300 0.000 775.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 746.260 0.000 749.800 1.120 ;
  LAYER metal3 ;
  RECT 746.260 0.000 749.800 1.120 ;
  LAYER metal2 ;
  RECT 746.260 0.000 749.800 1.120 ;
  LAYER metal1 ;
  RECT 746.260 0.000 749.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 729.520 0.000 733.060 1.120 ;
  LAYER metal3 ;
  RECT 729.520 0.000 733.060 1.120 ;
  LAYER metal2 ;
  RECT 729.520 0.000 733.060 1.120 ;
  LAYER metal1 ;
  RECT 729.520 0.000 733.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.860 0.000 706.400 1.120 ;
  LAYER metal3 ;
  RECT 702.860 0.000 706.400 1.120 ;
  LAYER metal2 ;
  RECT 702.860 0.000 706.400 1.120 ;
  LAYER metal1 ;
  RECT 702.860 0.000 706.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 681.160 0.000 684.700 1.120 ;
  LAYER metal3 ;
  RECT 681.160 0.000 684.700 1.120 ;
  LAYER metal2 ;
  RECT 681.160 0.000 684.700 1.120 ;
  LAYER metal1 ;
  RECT 681.160 0.000 684.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 568.320 0.000 571.860 1.120 ;
  LAYER metal3 ;
  RECT 568.320 0.000 571.860 1.120 ;
  LAYER metal2 ;
  RECT 568.320 0.000 571.860 1.120 ;
  LAYER metal1 ;
  RECT 568.320 0.000 571.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.620 0.000 550.160 1.120 ;
  LAYER metal3 ;
  RECT 546.620 0.000 550.160 1.120 ;
  LAYER metal2 ;
  RECT 546.620 0.000 550.160 1.120 ;
  LAYER metal1 ;
  RECT 546.620 0.000 550.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 519.340 0.000 522.880 1.120 ;
  LAYER metal3 ;
  RECT 519.340 0.000 522.880 1.120 ;
  LAYER metal2 ;
  RECT 519.340 0.000 522.880 1.120 ;
  LAYER metal1 ;
  RECT 519.340 0.000 522.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 510.660 0.000 514.200 1.120 ;
  LAYER metal3 ;
  RECT 510.660 0.000 514.200 1.120 ;
  LAYER metal2 ;
  RECT 510.660 0.000 514.200 1.120 ;
  LAYER metal1 ;
  RECT 510.660 0.000 514.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER metal3 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER metal2 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER metal1 ;
  RECT 482.760 0.000 486.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER metal3 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER metal2 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER metal1 ;
  RECT 465.400 0.000 468.940 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal3 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal2 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal1 ;
  RECT 366.200 0.000 369.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER metal3 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER metal2 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER metal1 ;
  RECT 318.460 0.000 322.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER metal1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 991.440 0.000 992.560 1.120 ;
  LAYER metal3 ;
  RECT 991.440 0.000 992.560 1.120 ;
  LAYER metal2 ;
  RECT 991.440 0.000 992.560 1.120 ;
  LAYER metal1 ;
  RECT 991.440 0.000 992.560 1.120 ;
 END
END DO63
PIN DI63
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 983.380 0.000 984.500 1.120 ;
  LAYER metal3 ;
  RECT 983.380 0.000 984.500 1.120 ;
  LAYER metal2 ;
  RECT 983.380 0.000 984.500 1.120 ;
  LAYER metal1 ;
  RECT 983.380 0.000 984.500 1.120 ;
 END
END DI63
PIN DO62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER metal3 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER metal2 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER metal1 ;
  RECT 978.420 0.000 979.540 1.120 ;
 END
END DO62
PIN DI62
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 969.740 0.000 970.860 1.120 ;
  LAYER metal3 ;
  RECT 969.740 0.000 970.860 1.120 ;
  LAYER metal2 ;
  RECT 969.740 0.000 970.860 1.120 ;
  LAYER metal1 ;
  RECT 969.740 0.000 970.860 1.120 ;
 END
END DI62
PIN DO61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 961.680 0.000 962.800 1.120 ;
  LAYER metal3 ;
  RECT 961.680 0.000 962.800 1.120 ;
  LAYER metal2 ;
  RECT 961.680 0.000 962.800 1.120 ;
  LAYER metal1 ;
  RECT 961.680 0.000 962.800 1.120 ;
 END
END DO61
PIN DI61
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 953.000 0.000 954.120 1.120 ;
  LAYER metal3 ;
  RECT 953.000 0.000 954.120 1.120 ;
  LAYER metal2 ;
  RECT 953.000 0.000 954.120 1.120 ;
  LAYER metal1 ;
  RECT 953.000 0.000 954.120 1.120 ;
 END
END DI61
PIN DO60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 948.040 0.000 949.160 1.120 ;
  LAYER metal3 ;
  RECT 948.040 0.000 949.160 1.120 ;
  LAYER metal2 ;
  RECT 948.040 0.000 949.160 1.120 ;
  LAYER metal1 ;
  RECT 948.040 0.000 949.160 1.120 ;
 END
END DO60
PIN DI60
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal3 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal2 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal1 ;
  RECT 939.980 0.000 941.100 1.120 ;
 END
END DI60
PIN DO59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 935.020 0.000 936.140 1.120 ;
  LAYER metal3 ;
  RECT 935.020 0.000 936.140 1.120 ;
  LAYER metal2 ;
  RECT 935.020 0.000 936.140 1.120 ;
  LAYER metal1 ;
  RECT 935.020 0.000 936.140 1.120 ;
 END
END DO59
PIN DI59
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 926.340 0.000 927.460 1.120 ;
  LAYER metal3 ;
  RECT 926.340 0.000 927.460 1.120 ;
  LAYER metal2 ;
  RECT 926.340 0.000 927.460 1.120 ;
  LAYER metal1 ;
  RECT 926.340 0.000 927.460 1.120 ;
 END
END DI59
PIN DO58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal3 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal2 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal1 ;
  RECT 922.000 0.000 923.120 1.120 ;
 END
END DO58
PIN DI58
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal3 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal2 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal1 ;
  RECT 913.320 0.000 914.440 1.120 ;
 END
END DI58
PIN DO57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 905.260 0.000 906.380 1.120 ;
  LAYER metal3 ;
  RECT 905.260 0.000 906.380 1.120 ;
  LAYER metal2 ;
  RECT 905.260 0.000 906.380 1.120 ;
  LAYER metal1 ;
  RECT 905.260 0.000 906.380 1.120 ;
 END
END DO57
PIN DI57
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 896.580 0.000 897.700 1.120 ;
  LAYER metal3 ;
  RECT 896.580 0.000 897.700 1.120 ;
  LAYER metal2 ;
  RECT 896.580 0.000 897.700 1.120 ;
  LAYER metal1 ;
  RECT 896.580 0.000 897.700 1.120 ;
 END
END DI57
PIN DO56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 891.620 0.000 892.740 1.120 ;
  LAYER metal3 ;
  RECT 891.620 0.000 892.740 1.120 ;
  LAYER metal2 ;
  RECT 891.620 0.000 892.740 1.120 ;
  LAYER metal1 ;
  RECT 891.620 0.000 892.740 1.120 ;
 END
END DO56
PIN DI56
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 883.560 0.000 884.680 1.120 ;
  LAYER metal3 ;
  RECT 883.560 0.000 884.680 1.120 ;
  LAYER metal2 ;
  RECT 883.560 0.000 884.680 1.120 ;
  LAYER metal1 ;
  RECT 883.560 0.000 884.680 1.120 ;
 END
END DI56
PIN DO55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 878.600 0.000 879.720 1.120 ;
  LAYER metal3 ;
  RECT 878.600 0.000 879.720 1.120 ;
  LAYER metal2 ;
  RECT 878.600 0.000 879.720 1.120 ;
  LAYER metal1 ;
  RECT 878.600 0.000 879.720 1.120 ;
 END
END DO55
PIN DI55
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 869.920 0.000 871.040 1.120 ;
  LAYER metal3 ;
  RECT 869.920 0.000 871.040 1.120 ;
  LAYER metal2 ;
  RECT 869.920 0.000 871.040 1.120 ;
  LAYER metal1 ;
  RECT 869.920 0.000 871.040 1.120 ;
 END
END DI55
PIN DO54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 864.960 0.000 866.080 1.120 ;
  LAYER metal3 ;
  RECT 864.960 0.000 866.080 1.120 ;
  LAYER metal2 ;
  RECT 864.960 0.000 866.080 1.120 ;
  LAYER metal1 ;
  RECT 864.960 0.000 866.080 1.120 ;
 END
END DO54
PIN DI54
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 856.900 0.000 858.020 1.120 ;
  LAYER metal3 ;
  RECT 856.900 0.000 858.020 1.120 ;
  LAYER metal2 ;
  RECT 856.900 0.000 858.020 1.120 ;
  LAYER metal1 ;
  RECT 856.900 0.000 858.020 1.120 ;
 END
END DI54
PIN DO53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 848.840 0.000 849.960 1.120 ;
  LAYER metal3 ;
  RECT 848.840 0.000 849.960 1.120 ;
  LAYER metal2 ;
  RECT 848.840 0.000 849.960 1.120 ;
  LAYER metal1 ;
  RECT 848.840 0.000 849.960 1.120 ;
 END
END DO53
PIN DI53
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 840.160 0.000 841.280 1.120 ;
  LAYER metal3 ;
  RECT 840.160 0.000 841.280 1.120 ;
  LAYER metal2 ;
  RECT 840.160 0.000 841.280 1.120 ;
  LAYER metal1 ;
  RECT 840.160 0.000 841.280 1.120 ;
 END
END DI53
PIN DO52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 835.200 0.000 836.320 1.120 ;
  LAYER metal3 ;
  RECT 835.200 0.000 836.320 1.120 ;
  LAYER metal2 ;
  RECT 835.200 0.000 836.320 1.120 ;
  LAYER metal1 ;
  RECT 835.200 0.000 836.320 1.120 ;
 END
END DO52
PIN DI52
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 827.140 0.000 828.260 1.120 ;
  LAYER metal3 ;
  RECT 827.140 0.000 828.260 1.120 ;
  LAYER metal2 ;
  RECT 827.140 0.000 828.260 1.120 ;
  LAYER metal1 ;
  RECT 827.140 0.000 828.260 1.120 ;
 END
END DI52
PIN DO51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 822.180 0.000 823.300 1.120 ;
  LAYER metal3 ;
  RECT 822.180 0.000 823.300 1.120 ;
  LAYER metal2 ;
  RECT 822.180 0.000 823.300 1.120 ;
  LAYER metal1 ;
  RECT 822.180 0.000 823.300 1.120 ;
 END
END DO51
PIN DI51
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 813.500 0.000 814.620 1.120 ;
  LAYER metal3 ;
  RECT 813.500 0.000 814.620 1.120 ;
  LAYER metal2 ;
  RECT 813.500 0.000 814.620 1.120 ;
  LAYER metal1 ;
  RECT 813.500 0.000 814.620 1.120 ;
 END
END DI51
PIN DO50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 808.540 0.000 809.660 1.120 ;
  LAYER metal3 ;
  RECT 808.540 0.000 809.660 1.120 ;
  LAYER metal2 ;
  RECT 808.540 0.000 809.660 1.120 ;
  LAYER metal1 ;
  RECT 808.540 0.000 809.660 1.120 ;
 END
END DO50
PIN DI50
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 800.480 0.000 801.600 1.120 ;
  LAYER metal3 ;
  RECT 800.480 0.000 801.600 1.120 ;
  LAYER metal2 ;
  RECT 800.480 0.000 801.600 1.120 ;
  LAYER metal1 ;
  RECT 800.480 0.000 801.600 1.120 ;
 END
END DI50
PIN DO49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 791.800 0.000 792.920 1.120 ;
  LAYER metal3 ;
  RECT 791.800 0.000 792.920 1.120 ;
  LAYER metal2 ;
  RECT 791.800 0.000 792.920 1.120 ;
  LAYER metal1 ;
  RECT 791.800 0.000 792.920 1.120 ;
 END
END DO49
PIN DI49
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 783.740 0.000 784.860 1.120 ;
  LAYER metal3 ;
  RECT 783.740 0.000 784.860 1.120 ;
  LAYER metal2 ;
  RECT 783.740 0.000 784.860 1.120 ;
  LAYER metal1 ;
  RECT 783.740 0.000 784.860 1.120 ;
 END
END DI49
PIN DO48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal3 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal2 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal1 ;
  RECT 778.780 0.000 779.900 1.120 ;
 END
END DO48
PIN DI48
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 770.100 0.000 771.220 1.120 ;
  LAYER metal3 ;
  RECT 770.100 0.000 771.220 1.120 ;
  LAYER metal2 ;
  RECT 770.100 0.000 771.220 1.120 ;
  LAYER metal1 ;
  RECT 770.100 0.000 771.220 1.120 ;
 END
END DI48
PIN DO47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 765.760 0.000 766.880 1.120 ;
  LAYER metal3 ;
  RECT 765.760 0.000 766.880 1.120 ;
  LAYER metal2 ;
  RECT 765.760 0.000 766.880 1.120 ;
  LAYER metal1 ;
  RECT 765.760 0.000 766.880 1.120 ;
 END
END DO47
PIN DI47
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 757.080 0.000 758.200 1.120 ;
  LAYER metal3 ;
  RECT 757.080 0.000 758.200 1.120 ;
  LAYER metal2 ;
  RECT 757.080 0.000 758.200 1.120 ;
  LAYER metal1 ;
  RECT 757.080 0.000 758.200 1.120 ;
 END
END DI47
PIN DO46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal3 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal2 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal1 ;
  RECT 752.120 0.000 753.240 1.120 ;
 END
END DO46
PIN DI46
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 744.060 0.000 745.180 1.120 ;
  LAYER metal3 ;
  RECT 744.060 0.000 745.180 1.120 ;
  LAYER metal2 ;
  RECT 744.060 0.000 745.180 1.120 ;
  LAYER metal1 ;
  RECT 744.060 0.000 745.180 1.120 ;
 END
END DI46
PIN DO45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 735.380 0.000 736.500 1.120 ;
  LAYER metal3 ;
  RECT 735.380 0.000 736.500 1.120 ;
  LAYER metal2 ;
  RECT 735.380 0.000 736.500 1.120 ;
  LAYER metal1 ;
  RECT 735.380 0.000 736.500 1.120 ;
 END
END DO45
PIN DI45
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 727.320 0.000 728.440 1.120 ;
  LAYER metal3 ;
  RECT 727.320 0.000 728.440 1.120 ;
  LAYER metal2 ;
  RECT 727.320 0.000 728.440 1.120 ;
  LAYER metal1 ;
  RECT 727.320 0.000 728.440 1.120 ;
 END
END DI45
PIN DO44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 722.360 0.000 723.480 1.120 ;
  LAYER metal3 ;
  RECT 722.360 0.000 723.480 1.120 ;
  LAYER metal2 ;
  RECT 722.360 0.000 723.480 1.120 ;
  LAYER metal1 ;
  RECT 722.360 0.000 723.480 1.120 ;
 END
END DO44
PIN DI44
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 713.680 0.000 714.800 1.120 ;
  LAYER metal3 ;
  RECT 713.680 0.000 714.800 1.120 ;
  LAYER metal2 ;
  RECT 713.680 0.000 714.800 1.120 ;
  LAYER metal1 ;
  RECT 713.680 0.000 714.800 1.120 ;
 END
END DI44
PIN DO43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 708.720 0.000 709.840 1.120 ;
  LAYER metal3 ;
  RECT 708.720 0.000 709.840 1.120 ;
  LAYER metal2 ;
  RECT 708.720 0.000 709.840 1.120 ;
  LAYER metal1 ;
  RECT 708.720 0.000 709.840 1.120 ;
 END
END DO43
PIN DI43
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 700.660 0.000 701.780 1.120 ;
  LAYER metal3 ;
  RECT 700.660 0.000 701.780 1.120 ;
  LAYER metal2 ;
  RECT 700.660 0.000 701.780 1.120 ;
  LAYER metal1 ;
  RECT 700.660 0.000 701.780 1.120 ;
 END
END DI43
PIN DO42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal3 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal2 ;
  RECT 695.700 0.000 696.820 1.120 ;
  LAYER metal1 ;
  RECT 695.700 0.000 696.820 1.120 ;
 END
END DO42
PIN DI42
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal3 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal2 ;
  RECT 687.020 0.000 688.140 1.120 ;
  LAYER metal1 ;
  RECT 687.020 0.000 688.140 1.120 ;
 END
END DI42
PIN DO41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 678.960 0.000 680.080 1.120 ;
  LAYER metal3 ;
  RECT 678.960 0.000 680.080 1.120 ;
  LAYER metal2 ;
  RECT 678.960 0.000 680.080 1.120 ;
  LAYER metal1 ;
  RECT 678.960 0.000 680.080 1.120 ;
 END
END DO41
PIN DI41
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 670.900 0.000 672.020 1.120 ;
  LAYER metal3 ;
  RECT 670.900 0.000 672.020 1.120 ;
  LAYER metal2 ;
  RECT 670.900 0.000 672.020 1.120 ;
  LAYER metal1 ;
  RECT 670.900 0.000 672.020 1.120 ;
 END
END DI41
PIN DO40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 665.940 0.000 667.060 1.120 ;
  LAYER metal3 ;
  RECT 665.940 0.000 667.060 1.120 ;
  LAYER metal2 ;
  RECT 665.940 0.000 667.060 1.120 ;
  LAYER metal1 ;
  RECT 665.940 0.000 667.060 1.120 ;
 END
END DO40
PIN DI40
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 657.260 0.000 658.380 1.120 ;
  LAYER metal3 ;
  RECT 657.260 0.000 658.380 1.120 ;
  LAYER metal2 ;
  RECT 657.260 0.000 658.380 1.120 ;
  LAYER metal1 ;
  RECT 657.260 0.000 658.380 1.120 ;
 END
END DI40
PIN DO39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal3 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal2 ;
  RECT 652.300 0.000 653.420 1.120 ;
  LAYER metal1 ;
  RECT 652.300 0.000 653.420 1.120 ;
 END
END DO39
PIN DI39
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal3 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal2 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal1 ;
  RECT 644.240 0.000 645.360 1.120 ;
 END
END DI39
PIN DO38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal3 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal2 ;
  RECT 639.280 0.000 640.400 1.120 ;
  LAYER metal1 ;
  RECT 639.280 0.000 640.400 1.120 ;
 END
END DO38
PIN DI38
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal3 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal2 ;
  RECT 630.600 0.000 631.720 1.120 ;
  LAYER metal1 ;
  RECT 630.600 0.000 631.720 1.120 ;
 END
END DI38
PIN DO37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 622.540 0.000 623.660 1.120 ;
  LAYER metal3 ;
  RECT 622.540 0.000 623.660 1.120 ;
  LAYER metal2 ;
  RECT 622.540 0.000 623.660 1.120 ;
  LAYER metal1 ;
  RECT 622.540 0.000 623.660 1.120 ;
 END
END DO37
PIN DI37
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER metal3 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER metal2 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER metal1 ;
  RECT 613.860 0.000 614.980 1.120 ;
 END
END DI37
PIN DO36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 608.900 0.000 610.020 1.120 ;
  LAYER metal3 ;
  RECT 608.900 0.000 610.020 1.120 ;
  LAYER metal2 ;
  RECT 608.900 0.000 610.020 1.120 ;
  LAYER metal1 ;
  RECT 608.900 0.000 610.020 1.120 ;
 END
END DO36
PIN DI36
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 600.840 0.000 601.960 1.120 ;
  LAYER metal3 ;
  RECT 600.840 0.000 601.960 1.120 ;
  LAYER metal2 ;
  RECT 600.840 0.000 601.960 1.120 ;
  LAYER metal1 ;
  RECT 600.840 0.000 601.960 1.120 ;
 END
END DI36
PIN DO35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal3 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal2 ;
  RECT 595.880 0.000 597.000 1.120 ;
  LAYER metal1 ;
  RECT 595.880 0.000 597.000 1.120 ;
 END
END DO35
PIN DI35
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal3 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal2 ;
  RECT 587.820 0.000 588.940 1.120 ;
  LAYER metal1 ;
  RECT 587.820 0.000 588.940 1.120 ;
 END
END DI35
PIN DO34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal3 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal2 ;
  RECT 582.860 0.000 583.980 1.120 ;
  LAYER metal1 ;
  RECT 582.860 0.000 583.980 1.120 ;
 END
END DO34
PIN DI34
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal3 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal2 ;
  RECT 574.180 0.000 575.300 1.120 ;
  LAYER metal1 ;
  RECT 574.180 0.000 575.300 1.120 ;
 END
END DI34
PIN DO33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 566.120 0.000 567.240 1.120 ;
  LAYER metal3 ;
  RECT 566.120 0.000 567.240 1.120 ;
  LAYER metal2 ;
  RECT 566.120 0.000 567.240 1.120 ;
  LAYER metal1 ;
  RECT 566.120 0.000 567.240 1.120 ;
 END
END DO33
PIN DI33
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal3 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal2 ;
  RECT 557.440 0.000 558.560 1.120 ;
  LAYER metal1 ;
  RECT 557.440 0.000 558.560 1.120 ;
 END
END DI33
PIN DO32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 552.480 0.000 553.600 1.120 ;
  LAYER metal3 ;
  RECT 552.480 0.000 553.600 1.120 ;
  LAYER metal2 ;
  RECT 552.480 0.000 553.600 1.120 ;
  LAYER metal1 ;
  RECT 552.480 0.000 553.600 1.120 ;
 END
END DO32
PIN DI32
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal3 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal2 ;
  RECT 544.420 0.000 545.540 1.120 ;
  LAYER metal1 ;
  RECT 544.420 0.000 545.540 1.120 ;
 END
END DI32
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER metal3 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER metal2 ;
  RECT 538.840 0.000 539.960 1.120 ;
  LAYER metal1 ;
  RECT 538.840 0.000 539.960 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal3 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal2 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal1 ;
  RECT 536.980 0.000 538.100 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 532.020 0.000 533.140 1.120 ;
  LAYER metal3 ;
  RECT 532.020 0.000 533.140 1.120 ;
  LAYER metal2 ;
  RECT 532.020 0.000 533.140 1.120 ;
  LAYER metal1 ;
  RECT 532.020 0.000 533.140 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 530.160 0.000 531.280 1.120 ;
  LAYER metal3 ;
  RECT 530.160 0.000 531.280 1.120 ;
  LAYER metal2 ;
  RECT 530.160 0.000 531.280 1.120 ;
  LAYER metal1 ;
  RECT 530.160 0.000 531.280 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 508.460 0.000 509.580 1.120 ;
  LAYER metal3 ;
  RECT 508.460 0.000 509.580 1.120 ;
  LAYER metal2 ;
  RECT 508.460 0.000 509.580 1.120 ;
  LAYER metal1 ;
  RECT 508.460 0.000 509.580 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 505.360 0.000 506.480 1.120 ;
  LAYER metal3 ;
  RECT 505.360 0.000 506.480 1.120 ;
  LAYER metal2 ;
  RECT 505.360 0.000 506.480 1.120 ;
  LAYER metal1 ;
  RECT 505.360 0.000 506.480 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 502.880 0.000 504.000 1.120 ;
  LAYER metal3 ;
  RECT 502.880 0.000 504.000 1.120 ;
  LAYER metal2 ;
  RECT 502.880 0.000 504.000 1.120 ;
  LAYER metal1 ;
  RECT 502.880 0.000 504.000 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER metal3 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER metal2 ;
  RECT 499.160 0.000 500.280 1.120 ;
  LAYER metal1 ;
  RECT 499.160 0.000 500.280 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal3 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal2 ;
  RECT 491.100 0.000 492.220 1.120 ;
  LAYER metal1 ;
  RECT 491.100 0.000 492.220 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER metal3 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER metal2 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER metal1 ;
  RECT 480.560 0.000 481.680 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER metal3 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER metal2 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER metal1 ;
  RECT 477.460 0.000 478.580 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER metal3 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER metal2 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER metal1 ;
  RECT 470.020 0.000 471.140 1.120 ;
 END
END A8
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER metal3 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER metal2 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER metal1 ;
  RECT 458.860 0.000 459.980 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER metal3 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER metal2 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER metal1 ;
  RECT 450.800 0.000 451.920 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER metal3 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER metal2 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER metal1 ;
  RECT 445.840 0.000 446.960 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER metal3 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER metal2 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER metal1 ;
  RECT 437.160 0.000 438.280 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER metal3 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER metal2 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER metal1 ;
  RECT 420.420 0.000 421.540 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER metal3 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER metal2 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER metal1 ;
  RECT 415.460 0.000 416.580 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER metal3 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER metal2 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER metal1 ;
  RECT 407.400 0.000 408.520 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER metal3 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER metal2 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER metal1 ;
  RECT 393.760 0.000 394.880 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER metal3 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER metal2 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER metal1 ;
  RECT 389.420 0.000 390.540 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER metal3 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER metal2 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER metal1 ;
  RECT 380.740 0.000 381.860 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal3 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal2 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal1 ;
  RECT 350.980 0.000 352.100 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER metal3 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER metal2 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER metal1 ;
  RECT 346.020 0.000 347.140 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal3 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal2 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal1 ;
  RECT 337.340 0.000 338.460 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER metal3 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER metal2 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER metal1 ;
  RECT 332.380 0.000 333.500 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER metal3 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER metal2 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER metal1 ;
  RECT 324.320 0.000 325.440 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal3 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal2 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal1 ;
  RECT 316.260 0.000 317.380 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER metal3 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER metal2 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER metal1 ;
  RECT 307.580 0.000 308.700 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal3 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal2 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER metal1 ;
  RECT 302.620 0.000 303.740 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal3 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal2 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER metal1 ;
  RECT 294.560 0.000 295.680 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER metal1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal3 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal2 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER metal1 ;
  RECT 280.920 0.000 282.040 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI16
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 1005.020 294.000 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 1005.020 294.000 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 1005.020 294.000 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 1005.020 294.000 ;
  LAYER via ;
  RECT 0.000 0.140 1005.020 294.000 ;
  LAYER via2 ;
  RECT 0.000 0.140 1005.020 294.000 ;
  LAYER via3 ;
  RECT 0.000 0.140 1005.020 294.000 ;
END
END SUMA180_512X64X1BM1
END LIBRARY



