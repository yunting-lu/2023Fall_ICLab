//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab04 Exercise		: Siamese Neural Network
//   Author     		: Jia-Yu Lee (maggie8905121@gmail.com)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2023-09)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME      70.0
`define SEED_NUMBER     28825252
`define PATTERN_NUMBER 100

module PATTERN(
    //Output Port
    clk,
    rst_n,
    //cg_en,
    in_valid,
    Img,
    Kernel,
	Weight,
    Opt,
    //Input Port
    out_valid,
    out
    );


`protected
+?-2]+ZN_G)L+e\YDF;SW;KFD/7.I3Sa2@XM;SaUea;Z3A&fHd[I.)6-;aT?RKgb
S3GZV=_Qb@d/#B_J&B_=([(;)TM[[,EZ7^ZE(79I9Y[CJJ4O/ALR3^UG;Of@+K[g
WM<PFdbe@>>c\22Z(0&)P>-Z=BPe<F>;B813MJ^Ag]A#)8XP7_1f2d.5>A(.+V]6
+AeP5(&M+]P1B3\<e)/ULc_AAPJSYaNY4OYHe^:P8Y/T>WS;(-fOM?FI2@f[^Q/d
eVF:)_<8^9@WgGR]bC-&-F_[07e\E0e5-9H8S_eAR9=#KU;<F:,^-dFIK$
`endprotected
output          clk, rst_n, in_valid;

`protected
[YfVd&R)_#_LRL;D(95E#4NNT/1#^@8-FF0Y7^SWgWc&eK><4aYQ))<)3UL4]0YZ
WNSd:UXYQ-(bKFf3-IRGfY]KVa(_R,VbKQ?2g00.cO6&F$
`endprotected
output  [31:0]  Img;
output  [31:0]  Kernel;
output  [31:0]  Weight;
output  [ 1:0]  Opt;
input           out_valid;
input   [31:0]  out;


`protected
\V^-0F?.;RC;dBIff19R.f2Dd+^5ZW0GQX\,<de\bV#\3F[:5TYS&);0_,CA8V@L
gX]C&NI=ZX/N_LTG1P_FVe^N)QA:0BT-;2W>eeE:?SDZCPIPB[H.M)fDg6C,)2:3
eKg)\@AX.=)Xa?Q5IIE.S@GGJe;FLE_?7(KPB=QNCE\EgV+Y4]K&ZV&Y=/-J2Ma[
N<<0OTOIKWS]CF1XY4:TWAU0<1^2JWY6+L^YfM]Y@DQUcb:c@9=FdM_7aT1@1W64
4ZK,^c+^VLQ&JSc;05PXLDfDF.:JfKOT,8X^3d36WET-Je,#,D0^>@[VEf?4Z#AR
OAIXXKg(Md4#IN8YGg:<9gRQ;02CQL/PgF,-aF0F-NQ&;S.GOSP3=@\AEf/2c^TZ
(CHE@Y2EE6-V(\?@-XYG65.#:KGU3S,UFM[3P<1c:IZ1Mad171e-EQ.94M&K;&)I
dP]2/P3-Jc;=-3Y]MX-RRVB5SU7I)Q:6=74]QO.U,W5d]NHN#QJJT;)ee\dN)/8M
7U@Bg>-ED.6QTf<5d<]Hf()&71;&D;)RQL:.[c.75]-?aT?J221Y-<d57Y-U1DXa
gTg>KKK?Z?8g1YZ;63-cKBH<;S#L:\.U&=]]eTROSV-6)ZQ]cB;4Q^>&5Y<1K.GO
T,#5VFdf5,X.U_K?=?0C:]_SMbcI?W<8JQc:O(35G.BY)E:2f;cKJ<\M)f)JU2.B
a5<3L,,Kge#<>\MeE9G\:6\76?Q\Gb<IR]b[I(e#^A?,\<CC6;WJdd[g7A18U36O
SQ:4bGXA6H_IV6LEIHVVWGeTAA/:=6W(d]bH2G]W?(2+_?_]1+I.WV0TSg;aS2c3
(+gN+P\6&DK]0SbJS5.&a0Q8V&dXE4H3F.7X7eCdWFX\AOW]AdJW^8]VaM+N1I=>
NSdY3ALOHX__7BaB9;O)E(W4J#._P(&2,I0-9Q_UAFE0(eMV6ZL5YT.=,X=KZN8G
#,ea4b_PKa8]-(+C+3#Hg0,GGY_Ig-N:e8#]QD&T+FZW0LLV.CD[M0)V@./8>3&N
>])6@&,[+ga<>P0SY-QC<CR\MEM+fbb\bKDCY1E6PDDEH/7/6D47J;T6&O;US&d+
2cP#:?M1@/:gK.<&9/@/+9TWbEaDdS22=I,Z_,Fd?C3-H8Ve/U?A-0?CCN1.Y._:
FVK?\4NOZT&VcdT7]),2Z9eRK2ONWF1^=Q4R3+?G79170?8B=]6g4BJ>ZAP.8DKH
KJLV8<YIYf@[M57@/387RVOIDY?HFGSN=GCXKgAXCL6&2S&7#7JYV-R8/\&DT4d-
g&G-6gMV9U>5_L]BZ\<295WaMTQM@b1]TE<Q/3,9S6:@&C_J;)^Z(D?JU]Q)4Qdb
IaJa(Y])&\DO-,0aV^Acc&]/SLZQc=BI2L)\?/7g:OUW6Na_Hcb)PaXJ3g+1c5V\
5VU8b9\9CC,QA4/\6Pg#7e[)-I,]aA<c&AN-JgV1d#XbBZW4Z(<4W;)7<?RZ[#)T
f2O3XNO>(,8TV>KS#f0dR:92YbX2N?;H6??9UA,K6RB+a<Q4D+#g(VAT8KI;BM4+
38Nb^22@1g-e[g_VbC]-8J2@@Yc5=?A_eJ[NF<7-IY;8UHM8YA_-<-6^F5;(GK;#
69[-NN+F<KL01-N&QYeeM7ON]SgM@UZPOHCFHWDF(Y>=FSK&;cG3B]MB_(D@;Tf1
NEM/6K58H0#S@Q1U\4J6K_[(bS,=Q.51IPI(;L8J(C7MBH>fO0&1LVP81aGb+@X(
;)NZAf&1;\0aFF2Yb0LE&8R=X9TFK3g7cP?8XP&Nag<I:Wa\GG09KY,SdK)J,DGb
0:=CJI;RRNP;2-AQ+UW-^UVSKaJM4K\#W>e70&g>7)_C#2E-6CB&J3\@_97.J_JO
A,RT\b#]\E;264@D\.;G6D-F&CWA_.Cb9gCNcM/cId8LAN48df[6/G.254,(<C?d
P&]bF3#:&?Y)@0R+FF)B85gZD5Ub3NAEe\N.8E4#A?.W6+G.?SQc;KW89eC71ea+
CE>J40<>.7P8<H^^H290;VLZf\GP&P;dg>FJ-\;J+J3gIA_-\ZXQgObC_d#,>5NA
_O0e3TaWDG#Q.a(#E\-#91:d6>SfbWALQ\8Tc<^bQ/3=UU=YZ=K8#<]H7LgB>/fT
+:S?8[B7?)EcUTBR-(N;:Se>,Y7W/TT/504Q(+C+4CU&S=UW5MNZbH>9FL>e<^[=
cV;Be?\.HAL:e?@F&F,R#Y^>B@Ke_8RW;MB2J=SQaaCZecPR#JSDHDaX=.\(5D1E
^bf:I;IF96M[EL-4B6#?PCC2#;//2P)#.e+e\^<3I\0.C\c=I\H(@TIWgNZf.6IG
E=]7P.[N_[,0P6TD77JH#b[>BK#=LaO:&eEa:e[<&97)Yg+;bYb<R4,Hb@\F>&5H
\CgZVX?.)fP@A93DXU8SXI\V[B4MU#aHf.g^BKTX2V)+&cQ-33AJ=,9=ZQ32a>RA
U=TWG1MSF/eaLPDa9IIQW5Rd/D\=LFRQ[3=_b7DDQWg2aG2f?fO0V=4f8Q[-,3F]
I>PBNZe+@JeI3\A7ZS-<\_^AXD.10U,;30TK<bDa<;/2)F?CA1),fJ9GUgZW<=UE
bT/[>&)K9W:@5C;QTe;0/=:-/30#f=V(52>50;D9@G.11e(\5#<1bYfS-W[VTJF0
2?T]g6BYUgJ3C2&1X_?/MW^O-A&FZ=g,a0SMbB-+O(WAU6c[/(QSgX0TTXCTX]HP
g[EJ&e)LL3Aa_K?eN+DJ([>#^>TPB(022dg=;U[e4.;dQ2YGb[cL9I=9#]PJ@E1J
b\c78;;<B@P@KaH&G;8AIf39ab[GY:/#;POT]X@>@5NYG8T?+RKgVQC^S9P#3-cb
VPTb0A#.=US/YQVDIZ?R,GGgO^0bI5R?bC?Z(c->)L7:ZB@Oe(bOg,V>&9:QM?^;
:fF#AceU?dC5T//^\AEH,cSNZI#b-\aLIVK?^?X5+9D^(0(J_UHV-JQ2K]AX@ZBY
:Z9c.cB0QKG+AF/=-e^>0D;61O&58);Dd:Ode7=F>>9FR[8]IL7b+,NYZcgDH-1.
8O3.E\KTfHB#8g@@@F@+MXW7;_1=I/\)T-CP^]L^e.ceRb;O+8bP4W864-M5M.d3
?S#c[\\EN87L.X^dBOd>]9#FMQ8.KBE[J(USD^USR3+NLBFINIK_KVbM9>UMFeQA
/8^eD0gQ.5AL&d;,Y_8Z2]Z16E7(MM\1STB]O#^VL1OSJ9ED1=9WXG\7EA.(^+OM
5S2-d8<#bb=E416D;#:I(5bH5:Q+R-RZ\RZ-d:baSFI2>8[>/XfgKPWgX(B&U<.Q
-d=I[5@C7a,=<c.])KM(Z=>HP2)TJ,W)J?[(g:RZdF9I98E_@O,^fWK)?2Z=.HBU
J@5:J7DJNIH38JRO^1FZ8&E0^.QO@^bg@\(M]0>LEB:#@>]J&[f@2DC9Le04W)?L
H4EWZP7eX=ZMW)JL+DLMA-P:=Ya.ED7.3IKX_eD8;)[8c9<6FSRE,J5gec<G&OdL
N\J_&-W:aAO]JfP\H6F9JF:Y?\gHQVNBT=T7P_GYeCU=b#B<70.D+?9^)Jc202A9
gW&VCK:@?<#(D5=:FN<PX]JJ7LG6PO3.ed70FWMJ#P#bX]=X19\A&bM/2=PMX5SU
KJ)V#5G7DC-I5HEgfXX+3,Vf05<C3WP-.g-G^[0S[R\_^<@@P;a[EH^DB@71ad@[
ZbO)^(XK;CW(W#4MHf4R^:LN.(b[DS1::d.@\25W5RgKM:BS:[fT7>0PB3)cHI<?
#16H4bLM8B9&L.>J?,(Y?a-7b_+g1F1Y8-](F6?NW[aV=I[&\(cZ^?cA-L1gRQC6
g8)ADO3\g=NF?.W1U..VZX4Y4Q4bQQ>RHRA_#MYAKM1MP@@aJ2@a0_0@7P;5(:TJ
^7,/^7<RM7]a]^J\SYH+G>(,X;cfOGZe0K]Y;gEFAf^Hb<+>gT_IHJT-\<If]ABL
#E=#)^D,Ka1,(]U-f&_Ld9N?(RgDM7-,aN#YaH8-S+PV>;?YT<JISNZ-8GSf[4G-
,>VEGg=#MdR#HR9+dY)=Bc7VbF]0b@X+5c#E(X1\8O1L>??N#5fF.K6F^>g4c:OP
]:e(C63K:EHUI:/-1bWW^1.G;,WeL>XBO_62cND.eKL#,@1F@(AXg+)5f,.#>@9R
YPca\f28CN,_7KVEC_IC&:ALJ?009B:PfX\#8B\bdR_We>:>XJ_Y.:N8#PTXe-#H
JS[J_82gOHc&EC0TT(J\6^(=BTLLPdQ_=]EYK0RSZ[gG[PVS,\<?aT<OgOPPBY(+
Fc?Yg2ZNaWC@^8KG4X[HFQH]EJ_KJY2eLZGW0]VGb\E8W;Y-I)=7,PfE]BJR#^/H
R=JZ5_DT/2>]-DJa+G6?KVII:S)4XA;4C=;W^6H(&YY,D\G00,8FFBHSUg9L#M9U
a^G&:WcYK)9TVc[[VXf_cbXHT5)a+9Y]NXV.^_I6R#Y/2T1C#TaBQ(#\TX9O8M(T
SIAL=0f=ePCW3_V8O1=GUeCCV]?#CJV\D6FC7T<B)=SXc[UWd3H).H0UNbSD++RX
E3_OZ+E?+0NN7bWQZ)/_N3_34WAUEdJgN5MaJ1O])V@)VS]RTY&Ec6]R\#+1=dJ6
Bd=N0-4[fE:7B#9JAIB_73Ncb4TK4:c)>B))QReZ7@.L(gP_dQde7:1>BeMc3;>)
.H-f3:SV4=3W^2Jd(LJWe13dgMI8=R9FK0ZHWfQKV-^.-/9#06KR&&WL^_72a-CN
N9+FM+2Z&#XFTUI,_4If3?)V&aCScAC[>TPg1;-MRLLYI(TLc))@>I+A/<M]_4O+
73M[U#:Xc?\UI,:/d(I?OZ/^E8JIU;fd0M26U(^X]c<Hg?/76)6,RFfHS.Ld):V]
U=C?NdJM;1Z4NZY[]^ffI;Vd@]#&Kd4.\C7[JE^JVe61\P79T<G9E&)Zd5NTSP?Z
e&U8^N,e1eb87d=:0(;ZLDEH&_<7VYGJEC#JQ]<03aLU@1SU[Qa,)L]J+BC&C@58
<&TR9#[+:V[05].(N9]XWHaI)60:0&#,fTCA:e5B<65BF;F@H>S>_1bX/NLA@c<T
IG0NVGGbf@:VQf2/1Y>-F@R7D17WgfH1aVN^#4_)YC,6@+RZfMI<c0ZGdU?fN1aa
L;I36b#7D)(M[b-Lc5C6:aP@8g(Iaf8;5La7NDWb=)>TO)[1L&C)<0a;,9(?P+9Z
&O1b_Wb8facRRZ[8T/gMSR=.BF4;WG+56@-De5:U?HaZa46S&VEV@-cDO;L&M9d]
J2#KXF[W.^8DT15GeP<-M(#Q2&Sa?Z#57PLNLHBd],d<B;(I<F&D^g)V4)NSL2((
CGADY5[N)d=[H,9MP6ae-:]+0E:[^)USY;&gc,6>[F0;+3TW,&QfNG-2V+e<aH<X
1ge8MVfAbf:35FAS[^-Dg)#Yb=JSLT)NK]I;O#@2>f,DK69K9,1U]U=LTMX)4NMD
B/_F_Z^KXc8]a<Fd-9/JFf..,061J@J@2QFNSF[Hd1<L0PQ@M4D/UW;4Q4\UEf2d
dd&4(=1+Y,V+Dd;-?Bde#Y2fF#27c#fI4E[N\H\8FM,,g-HH2SaTONMKT?2c:Ta:
EVOQ3dWBMRX;9_\^=d\9M9XK46Y.VQd+.P<)9;8=4)3cS:\GAS1;]BeK,3SRO6T[
:GKY.fb.J1-Y\2cNN(QV\U.R31V7MHabS-7Wb9NG&JAXBHYYA@._IMaS#eQf;1:f
Q97VL0/fc<:0C/8][/#3>_Z0CV[41VP4Neg:aO)PZR,SYRRFIeJc5I1<M73(VPRH
S.62Y=CI.2B(N41MUQT)?]1A/G8^J<fAFD+d7-#.),)\KT^VIdCK#b[E6\fQRQ+^
2,FV[MM7^I[5V#=6/+0?\?UWFdDa.8BZTcU7a.+g\[EPaIC4f<RS)([dA8ZMFg33
EMTUUgVK26_=:Ege5G_K\[EJ.A8Q<4UUfM6f;A<TbZ2M-Y#;+E_^8:eINQGV^ZF8
I:7PUI#J-7QKT@4U]>gX;-I:N[C,RQ2O(QD,,JQEc>D0EW]Pf(9CcG[_=R>EJDRM
55FE+3#WPQ^IV=,84X]=4g+Jg^]+VgKA(1TMg?89]D)V-^KT7B?LgSKTDM[29K;<
8HD+-^dVO\^=0Ld)_U<IE4U/QS-7FVN1BS=8;LXKVQ3)d]/X.dagQZ?)OF1caZO+
-#S;0FGN:bDZGTb2C8SG=++PFgI?f2caJC)1L=Z8c]ZIf9WW^fZ>Ca<>38R4M1CJ
NFFC]\fA1@]9G?-@:[_@C,\QY?-_SRfQ+8=PGR:].0(BEf[eD;b?AH1@#[fb)XCc
@_Ig+7:FdOA.J(UcN>(4c.Z^F228>R)Q;O,XcYF^4-HJg=VR^JaaG_@]@MIT#CFc
7aP^659:J1#7A3I)XW[/S[=W]DL2@?&V1@)#-0>,13BB(.ZAYX]KB5@L@.?J>63F
TFUJER[0T;M2Sa/.e(R5P<O^LHd&3,f&WGC(:O6#P?A?<7?SER)>)IY+Pf-Y(,T6
Xc\01V.X;gaFd;K^5EPH&<R[/ZS3Z#6R&_#P]>I/L-K#OLK#4=N<6J8P6]#ISb_@
>)1BC(<<GY/VV#-=>S>9)6&RY9K-)a^#8XEe0DR^NMJSFDWV8Y?;&B4Bd9A526bQ
T&@G5a.J),AHg3[gd5M=VH#:K17TUX]eFN(<_gV9F>PJ9O]b=3[@Sd/F57?Y?SBF
,?G-KI,SN_JVYJ&GcLNBg[fK/#\8HfV@JC[+P+;<M.d>_G_G&OR-U7GgR=L4441K
VQ=8=/Y8ae<_/eRWKI]8K0ga0(+(TgS44a3NFHHG)dURF6g^/d3V=M=f.MgK9N14
UJRAE.^U?Uf>,4Le_/T@e-e]aC89,3IPRW2>fF7)aB.:R512M47X3CF]+U;IM^dA
V,-bNaLUFaZDI,=F39-Va)VZ@BW)7JXT#f>6GQ4OC869_U1?_C&&F.:ID<OYe20>
Da2_Y#0(UT)U7;@IDJMGFcR3HI(]CO]_@I^<#-4bGXK_Eg16[OfM#DDXaT_P^6;8
?VSV[L+#3J]D:]_3cW:RVI[0@.R[K#>&350.^JeQ4(YX1\49BEAJL;O#D)CZY64G
T8?FG)VK(:c>@8L,YI,):+36@3e6KO;BG#1YQN^,MZe5_[E2<PdA::RRgH+GI3UI
P0?0,-Oe:0FP/8d9fa5<NI@C+BN43?LK5-72CYXd+G8VD2KWA;\)LI9-8fPV&4c]
<ST_31BJKY?A:g1]<^S4TI(3bFKCEIC1RZ^8K0_R.CCB804NTLDB9Lc_U=-W_\5/
6/cYS4)K3+=JKWZL,-eYN>7e0YPSc:GY-XXd8^D/CfK4(N[\^_;0G-a47]V<08C4
<A=E/G.]8?[+?[&)Y6_4L_WS_/aKC(JP@(gW&FJ<LQ8-?CafW)g,(PP_S66..)T3
>G7E_J?Wc5W_d?O0N#=R^W#QL2CKKT5SEA9#(UDJL(\Ib6.FR>1M>52?@Y7f8B(T
A4P@W\M3@BB9>Hc7,HcXUGGG+;+][<VEY/O>>3[E<0Y1,cd/X;J+E^+F;45WbbIQ
ZT39NZe@O-EVAX]HA]IRLeIdfUEA1QLGAH5Ic9WDF\<A>bUa<.](6G3O[cf,2\KW
]&SBE79UK3=70[793d#N?Q:GZPe/+@+cbU>Q_dMQ-&eJPCCF-fUC::7ZKW-:Q&X_
)U&W;OMC>dN-E&Q(SCPCQcD=(3b7F3#SL5S6ceQ\B&:c0_:ZM7a&9U1VU/c\6#T+
MA/<4)OQaW>QVZD;E(f6;)(eB)E\JJOC)?g\VI0C&_#Vf.K,K,==WDO7HPYad#\7
@1.)4bad<\e-C@\dASUe4,gW?9)F.cT5\Z]&414MK2=M+Y8YQY[1XT?4A_E21KZ.
D1)Y+@1,V\R4UN9V(^PeVd5(;72P4BB_)&Y:IN2[H=\90d-60T04NB<QU41@b1O>
S_EF5><f9NETPJ\/DCU9\,F1G1O<^5K?AeT)E\:eP_0=FK:a_USU\J8M;OADGT[W
8)fS.OE0V.ZEbLK-/&C\_,X9STM\MC5;N-:CE2/S/02S^f,K)LL[51Z;B-;).G96
IP_Gb@.=0:MDI5TNMO3GW7O=>[H#7dQ)7LPG^1Z7gS72RTUd=S(KSVHfB71+)-D.
G4[6Z7EM:D;COU.RIXP<=RCTAdc&5#@f7bWT:cG#D/7]de&e>f^WJ)NTD&?JJg)]
44g>X^gd2#YKbFS+^f\E<-XVPOYOP4@1JH:9@1Ga4C-.4PNN#H3+bcDbIZ1);(bU
(4bZ:2855d4:T(SWe5RaVf3#(ScdgVPe2c(75fJ+(]8S)d7fC/[N]7BWI1JY--KW
>Lf9UN5a&[/a;P=:T0Y4fRHGL4e-TT;R3Fb8Nc^@L1_^U]gdI66EESb13@Od4GEY
_SH-b#3X<f#=[XJY/B:,(d&X0XfUBc_<\-AG0C7fD.Y(aYWe][1Xe/7fYa?f)5MF
/eO)?(JC6>7F05LDIgVB9f17A((9X+V-^SWHW[c>BHDB:DH7+3@T\0->6\[)E<HB
SV=456ZLO-EBE)6=acMRaEG3EM4<c/F+RVY]<0[VC,&1b=H)^4O;b8ZgJ9TS3F\d
c^W_0[7=],K?T-L#dcRKHKaD_Z@.3,@9I)K3==c(JT,+A3:9g:f\ZKGB=#Z8IOMU
)FL:HX\d,K[J]_.Mb3=&Ud>5_7Y#5YC@4LaC.5b5JAEbDBL&75>,L#OXHL/(O(3<
2dB@0?R=QUA890<f]CB_Q0#^eSG/e:HR=450//AFWZ3<eb6\3XV5D6&DR]Qf/91C
D6c,B_EU0F^JXIJZCRD-DCTWPH[edS1D_?\-<SKVL2>ZB5-_S3?K]\1Y\=DKb2[N
+3L</I/?IL.&HKMN#B>W-(E2=]/aB0WVX6A)BDH+[[b2D1b/PEZTg^LO+U=X@EF;
(?@b,f+M9;1@5K-,M;DL/;:<KI,&[28b(,62XBafV/PcOX[]R+,dbZI5-]EY_7#?
J_LY2NIE]T/2Fa2<U,NOf^M?^CM+AfUH#&EES23@J?/];(/\1AQU+e/_b.[B97(V
+Ab.T&6cW.[4X?+J\c>X00@?d6Cf#3?K,BI-f6KgA\d&7]SH4_cE?6<RIV,[?5De
S?c:WH@-:QNV1>QbA_S_H=,?E;)XC_M6?f<gY5X8(b5e1e.ZOF6)9>;V)ZcZ][&^
fg-cYS,F75R6G[MJ;@6X<aGbE]M.fZb(7_YA0g\cc7);C-F<a46UIU+<6=//JSX<
>^&S&;.0]9:SPQ;YedN4JA3\UW3-A0GN\FAQ6cHg:,UVeQT.MA+C2_29&H^5N9M)
7FF7U8YFW,S7]4WL@C;PLCJ(E[7&U#UCI9I55(VOGVJ>13[UcQHP>]]a5AL]]_YP
;dbF5YAQ7#;:X+>-B44#BR6X;G,AOY0+HN^#\5K>egePI7:f(<?IG&IWQS[_?^Fc
5AKG5D;).[Tc]>.Cc5:e5=)F.K-.69J3Z@T[1GE;O-3,\5Q^#AIV.fD>Y7d>9ddT
dJf^cU5V6[A4(a@^Ze+YDVS5RKO^a3a/G&:d:.3CPS:D:>Y\(_9^B]3-f2H52JXI
gJUNZcDBCTT>+E7#eGCOQ1#49SO1@2IV4.>60\Z[_P7RcAcRD+Zb.dbWe.H.&Td:
.1,,WOE,ca+Tfbc<,8T<8K,E3^\HQ,2AZc^D[D[[e+L-S@1\A#UJS^?@>f0D8_?)
SK0XH0-?.-4I=gZ7dc<NWZS@(cREW?P<e.8;OefB/fG_1G0dXON6fL0=Q#M:d_;A
8]6?cUMK\T]#=6Q+?Z49f4c7-XHAD[[c?PF+B2V=4N_5e#MJQV@_b.3BT6\99Yg(
c#aNM]SbT:FAe:3A/S6YIFce;E0F:;,2-/-7aS>5>X.?JK#2UX.;>ZR]8X)^29AD
(Hg<L7f-=e5QD^J6-AE@B8KP?>7Ee15LBMB9D>e=eP/E4^N>g#a+;\BD<eHIU.N,
]HM&42P/UK-1AG?;VXOO9I.,W;TC^JZ8[[1,1b=?cWXR(6SZ\@^ET381T6ULIL4P
2002^gP@H]G+Ae&[,Df:>Q:dJP>M)(d?F-QVIG6cQ>HTgb1)S&.aGF^W.1I7G:>^
T1ee#10ef>-0H1974LGE)5Z(#\:(N]+FOa/X;Ca>,>ff9QNaRfU-Gc6OE?)aB]W.
IA=2IHI[0VB(7Y1,DX0YKD1fC@1(P#DSJfJKMQC\:&^^4eUQG)ZbSNL-+Cdf[T;S
d9=,:(#J76,G)#2WaH4R71I.fIB6U53IA-VT8K>R?DO:aY(H:VY9:;bC7&E-5_+M
_REg>bR[&U>T?aJ]0G@9aZ5PF58@M3;7UP35&>G0&D)N=4G],g7CLU6,;SH@Of>g
@]f93e:F;gd=##C-/G+HMa+R?Y@;<_FL@^?.>QE4f:7:e+1&#L:6(Vf_B3Df+<GS
5\Qg?Y3UP5IUgLPN<@S,-I&^LS):(fC/EG&M,I@;9bAG>P@B,I0GG/(VD7aU]B3c
EEHPX/P;e)@Zc4>VeJVY.e,K0-GH:dQQ8WKGZW7N_F\U@GbaVc>?WG4(D/S(6RbV
A2/=]JfLEWe]c,D4K=a[(NIPdC,#d8=aLH(\U\MWX[3FIbQ<_>TBUW5U0RR)\e-K
Q#;DR=E2g:CO/5\,;>AR0T##@B-_f77=+7K;)^]5T4Z1O_?KAcDdV?R=P&BSV.;S
fPfZ-980];V+S=H6dF1G=SI]&5eZd2(&Jg73(+\>S<Q&Q0XE;;aY1W2;ISH?ZVdP
V/0(#IgLM^,befZW0D9gSLK9R8[\5SE[N-0-<^<[;1D=T;EIS^(A:e\#:MT479X\
Q&WY(@^PH[O1LRA,5dXd-a;g?R55R+PfE1_V4G/(VIAMWf_>Y<EeJff0cac5HcC#
HT=BS6E3>5V#<M]/S,D,?e;9IE_W?gOPG@IAeIW-bg)c-5,YIfba/@W2(eNe[UH0
)M^X=c\[T[\R.#gI+M1>\(9)6;(&gcQcbY_PfX-c^_NGJa;AN=fCB?)2X74J_3C<
a\MLT-D_-EaF9USQB:==>K5X@dZ[1B9J);Rc:CTA/&Q1>b+K=#5GB;/6#fIQ),\a
@F?J<;E[\+B#^;[BFbK,gB)09&W1@6<K#ZC8\V5\(M<<NGS@N(bW?94&;e&\6(=Q
5_Ie<7=6H;32#5P])>#<Zcc9S4DZZT-T=^WM..b9:4@PYG=]8](R::-=J]J;bY&f
f4J&+ZM2fTCQ4afTe6[/>.d3gIb9S^F/eM,3M4aA&]8&b&aT#^CU<Q(L[<4JeK[3
N(/&LN)gQf4_>8V]<Ae=3P.K>;[HDd@g+8TbM5G;5LUF9[/F+[=SN;;(@dR1+CV1
C8TDCNP>\S2AaUVWcJXO&12L>]/I91MCMa:(S4]:7^Z)@[;bb,ZW3>HUfgY2R[E]
7RWI]bW<R4NJ7MK3H?EZ34)W6>+JH2(#;Pb)G-JF,+4XgbY,9f//830>EI^_2KV+
SO44K+LLPJ+B^0a/TQg1CDSd?P5@3fEDAE#E1=Uf1-Z4UY]5E>bZHE)NQ9.gbB0Y
CQP42H5aaH@22CLe9=I9_/I:BQ3JV=+U-4AT0<)FM36G8SRX8VV]N->=:eY51=[N
3/J0c2D+[Wc#>:cB_S@_Z2#@)63G)S6C1f3S.[77-FW3RP^HW_MbRGE_bZJ-3_^X
fa-bTS0T>V7]c=a/0>HABgSA6][]W;,B?9dH4[)bf4HcKBC5L(H.RW:3D-E-1K9B
P<W-P]:GK:WN=5NLKSOdP9]\?cH>(H]WcXD7F5??&)??[[BcFT6^+;f^,OWM0<<R
8MH6J;68C7OJ]CXSRN@K@+;0/d[/d(8-(H?T/X];XeP][F1C3bT&)&E+XgR9LMKE
acO3c]U;UF#83V.Y;9G,WI1R3.6\a7R[_-fZ=V,_PLXe3UAVYV_UL:.WA\9gV[?X
^A&@b?.W>57+1R#_@N&J4M]:3:A[g-]LHF?(7[RD6=T@(8](?,5U[=<bb])cG>I\
DU;Z)Q9XTL)3Sc6T4;FSa/)\RS^6-1T>CGSZEH4@(@.g;7T3)d&S_.PN8cOP:BA1
+SOM>V-/KZBAZ,a]>g2.P0^8\I&Af9dEZI?=cNL.b]=(F7b3WY9AOAD^;6YO1a4c
TgeSUOTQaOdcD(A+UMK]JT@GUO_4DDY3=/S;7CM\)a]+Y@dX\]J(aQ^THUX_9GGE
MEFKC&BW@X[SA]_G;3RI3=eJUM)7a<_]cIM^gYL4.C9[WTeKa?R2;O<U2\8]T-c:
[8_)==QKD=59IOI#:[R3gU:gd)6U9]Pd;H55f5;U[L]CA360RS-YHCGfXM41dP>G
:Y.fM+Bf&V_+fY];C^LUI#=>E+Eef5F\LG5T7C?3Y@:H_b19/R,-M4,<4Nf1B(W?
I^#/;.7F-]MSg)I;e9(DL)[-5T1?YW];<e6:2AG8I[^K#;GIHcTFa,;d6OJgT5_J
S5c.:\8I&U14Y@CXOG-g^C9;+2M.OOEYHXV7G^6/JfCDD];9_:DRa5<;UZU)(Pg/
.OG,#Md(:a_H[QZ>#Xe30Q6R.4M39Md.E5f;g6O9_Ff3Tg78f:KbE@0E2aRU)0<:
Rd]4O&BGTCL4Y]e_<[:1?>Hd5+MY2>Pc,CLR32RH2;G9-4/)cU.(LU\ZB)Z]#c:J
d;]GF/.^5I<W9aQ+5+68PDU^N,9MTV.P5eQ6AI).IB1#SM,A]46)6&23SP44OR:O
ZZ7_>\5>RL>E]33DE4^UR^I;JI\.\NfQ/Z0MYOFA44e\/RG[V7(3;>ZTVb,E>KEK
WL596L1L1S6,2C;eaSE+#AJfO1IIe_R3e@L[<VNU[Hf)MGf>Q7:bPGK2+URD(T:Q
<<VO\^/J2V4A\P#ORNGgR]aK]@D<^bUF7W;H7WFf/+,RCB)2+SB.:W]E;>2<?J/M
F3(fDG[OE84]/Xa<;(8TQ+5AT[-(@cB&Rg/CQ1]77FL6<aQO.2bL^>49cBcF2?4X
NUZ<YAV)BTeG3c-&#aRXJNT_T10.)T(U0)<[C@ffAaf?^@cB[Pd\.&1LCPLM=-9]
a+WY4]P#.#Z&K[:G#&)@)_WF/cHPMAA<BM9XTOSNdKgQ1g0,e2FcFM#XY@0WI\,O
)^ASHVE(-&I_/6^[KP0T#Yfg/8J+,)WQCYY-^LZK:]D=SJ.c;g-6ERY<DBJ&8]>[
(V,J=O-JUD(G45/,3H:YbgE92A.0GG&YB_2[NNR;([(B=5<&,D054=N3<b)^b&I_
W6b_@0=NT#78dTAY=&=B&O)@fPV#Y26KPUK2U]AZ0_UZ,-+KGJ&cQN<eQ^SNH\?4
,-;G@H(;YS4].A;Y3]f#7KB0PObAf>CM1;F05c8&^C)9E\D9^e?4^+?I/T)/G5K3
SHMG<8[V(S?S?b-c9;/bY>7V=#.3?O?/=aXe@HZ<AD+5Gd0c,.>#72HSK<U6f?U/
<YY^VP8_-b8_+:0[JU0C9Ndf1<4QbB-XC@S>933K.W,g9Wc)QL2[G5Ega:/YSZ#>
(BFKW&^I9.H&\T[K^9OQE&4>P[Ue_]gcTCNE@=).N8g?<W2#U0Nf>,/bNU82>HV7
966;+ILK2Z3.X0<@8H;^4W#dNXF@^D:M1gY@>c;;OO4UPA2ZI>0N>M7Fa:E^[ZE^
UK63CC;]7B@D,4d#TM=?_QG[:7QDM;PP,T:/)_c@.C&+O3K\(X)0d]3<4:A>7\M_
=K#-e6REY[MKe5d\-=PK#DOFI,45a/IUL0QE<8\T[4BRSDS=7FKA:HY/21U(AcGb
-7?HJOT:Ua]P;VR0#TU0V@VV&Me7([G1>BFb.YOXRB7.T1NQd8g/5EBAMWMUfRS#
\)V\>]O8IL2<U[IYf,WY.?Rcb,PAM)FGAU+D\Td3Ba@6R+bF+NCO0E;MDADC=XHC
d?e@A,PRbHfD9W;McD?;1ET#:NUWMgdMX]]INB<XC)dXb\N36(D>X8S99cZ4S+[X
-4/ACJOe)8[.dMPPgP:L>S=]1(0XHUd,J<5<EgJ,c]cL[1NB(\QJ3@@^7?].W39N
/NU5_W[-)A?AKeQYEVI3:=B,9NT?K(]DAMQ55CB.:/1Z:7aD>62/I,^<E]Cb3YN_
[30c0Y52_W]?=IfgDM5=_S@g=WG#-@_QEYB.NQ:cTaC/,GX>#E&eWPSFK5>7>VI/
Z:EO<N:OURJSWc)LT.\^g>bH:5M#\KI[Hd\.0]PQ6U)KQCBYee,]?0[fXE5BHe.Y
_5L4D=,2NbB;R((R70UbR?.RcD;R/Abb0HADOgJ4DD[&53VFK(eICbJ36E#&>PEZ
fT^G;Z&KLBI0=6DKJ=LMNaULKX)D\CWR[WB99D00&@Y+TL6?2M2K@c[P2eZ:g-FF
bT[+G1@M@dO9<+S0^=A6^=O46M\A<9/>^LX<8_PWEBQB)84?A\YXRcD;KGMISKN5
]#cP]TFR,4B9G?2g]?4HR+UL@@,2SXVDBFHR._Y_T]:2YMTBMb;]O<b?##KI[aI:
/-69/.RZ&UX)N9>#Rg6^T@,,@)dV_)b,WDHHf&6Z3]3C=EdcIb)DT&_U.;:ME86(
L\Cd+.>#RZEXK#J;>V;/,GPgK5&[(]O<.N[CeAL>)d6PN1Ze\eA#V]?L3cI+4PD5
EMAL/=1Rg)WG4_A0GTdQ7;Z992GMS]5IC_TB>K2+CI1F3E+32N1cD1+3?cE>^T39
3<NO?7gX1L+c1aR@=]2QP4K>TU#Q;eV5JNYBE-B>M/cN3DW@;UX+];,M3>T_aI<a
-#O,.WeDT7M43Ce.KHK.\,Z^16O9S&8G4EF-[F=OA9^0Yab=#VC?SJ?(PX?TW-Q3
g7a>0BP,Eb?PWFUaagg[QUIS04+7]9U9T-<HG&d?;VA]5S0P:c1#;c_YA>Q&QMeY
;#&D<;2d3KYL:G;b\Vg=LZ?1FgAJ11(WE]8__5,MWL1+E8C9cB]^>\?^dMdEV^EQ
75&CEU],X41)\ZA+NST/QZRfeWU,&Bb\bfA=?<b&0)BeYVcO;_bC(M,&@Z3<47^E
TA(XME83LR\\ZNABNg9d5/X5Kc+7-.Uf0,3Y@K>.?#MVYU.2O9>2A6Q=AIH@,6A1
PX1&I>PH-<UUU=Q[7ZG:BQS^1;N+c27&SK=-X7BV#_;FKdN03K:fF2D&TG;S+\KZ
K.K3\(?@YX\<EdaQJdL:L\&#PZZU\Bd5AXc7V+]61R#C&2#[4==5YHNJFS8f\F);
,4A54V)bbd_ZDg:QPg+df=9A-+)TP,FCQ/B>>,ecKKVXREA?Q#8KAZ\L=&1]Yc(S
X97BMP8_KJ<GR\R@O@V2>eODf1K>ZDK_@X#a^92N-CI+_J[C\?10RbB_bQQXAZGY
SG3C7H:\DLS+1U?:WSC]16=,3gFfN]EZ5-VQ>F#fP&I,gfE[:EaeMbIP0+5@=<+M
5EP,4]0c/aMLI]=80dQA:cDW9D0RZ-&FVTacB)7WdTZLDUcJ237D)8+R9WLC-b/b
CMO/RdRDTPL2N4TK2I=fJ[4>V0B3@SWFG9>UXQeSe6WU<NYMB&C/]bL50LFZH?Yb
gG@QL^YF@NY@bDKO@TRID])P^K#Kd:a83\P8TP;8082A\ZA7+^[T=f)fC2:Y.&6P
.3.N/bJR9CT?:>7,3<+UA+&I1U:DZFW,C?W.^Z_#K12J&f\5^.DP)8Y-4-G5XHM+
RY/V@)P,0dfJB>0Ld3XIaZ_J1-Z:BQS8-g#U&,/+P8O?LOa]64BXH^afUd>6BG87
8S.]6I+P[cP7Y7[.9agbPWASGOR+T/]H->&]+?.TDdOFLKf<+ZX)\OBVWcb,7QP[
Ja_&HH:e<fGEU>NM/FgeWRDQA9_RN/K-&E5d?K\Vg/Fc:9?T8LX>^f^;GIMAd)FK
U?f6J\,0H/=#R=N;ZgAbH/@-M)XbZ_@P/IPO-7ce[J>b^C<Y/ZGZ9Y3fZU.aESd9
I\XI_)6A].D0S-\KL02^T[F,6.9M\e<d+_HB^P]^dS?^^?&MLX(3ZIGKC45,,IK\
g]B8^-.g>=:Z]B,V2D^YgBRGG=)6eGfASg9V(W4SY83M=/NGA:SfISX<2EV888DI
Ca(:XQ2C:M5eCK_FK62:e)EG<_OA?-[&&5g20I5?:6_JN2DQWY429N/UDSG>5WVa
8>G_8d>WMALGObb.180fWLg3K(#6O3bc1SOX&OVLJ.a/+#\;3IEH,d;,bFV?+2D(
##&:G+LRL6_-TNO\E9AHJ)E@I)BI,@XfX],Q>:TebH<5FN+IQHPWQ@-fd7?EWIDP
O@e_bb)E>bID?#ZaV[P:0e2@ZB2YX9cR@4JBDBJd_f3Ef4389fLQJfH(G.K5HC^<
CA+>^E,)?7=&2BcK.f910,K;G]RbCGE]23JY+a+UHXC-#MO16&dS.^>2]Z1NCQ/S
PD;E-8,O?9@f5RH,::XH=H&1L2WTK[<A=_f(]:7@0@6W6I_O\2c43Y/&YaO1@[VR
,<S_8QMLCeOFB#LWCAf1d@@J&RC6MUV#^Xaea6(BT/3?J]\MJc[W3E3<DG)7WH?\
J,0=8?aOdd_\ZfBPAOA8W+KY<cYG=eRYI+=9DOFX14e7Z<J6XIX[KCaH:I4ePD]E
.5@O;Od&37O35b0QYAH=:TDMS3XMb2A1?URFad\=7AAdd0M7_2T>[D;4O)NJU-QF
6-<c@N1]&VMYU51S2LRR7f\O93MH<RV]C[RV\FO6LT^eP>(SUQPM:F7^&.c7,J46
[gGaLQ7e-36X.ZLZRdC?^I<E10Lb9cOa[Xg>4NOXYd(Wd/9<R>G27f4b#]MIY?EX
F>I=0+V(JaKAgF=R3PFGIR.4f(/-A?GX^CQeMd8g5^3<XI>?BFH+1;5[0J2KP@G:
]W7B:[SKS2f3A_9-3d&?SYb9SVR?gK@0;gEg4K&/2IO@QL=X,P.[J2BY:>XPI:EN
(]CR=<)\E1N&(#EMPV[ef_Ab:9F9IbBB4VT/TdeN77\03VRfbZB?@V0=PU:SEG3+
I^QLM/>9a>O4bUbC#UdAZ(bF:N,ga.4SF.e\92C]>F\97(\71</57QG(X,g]>P]L
eKA78b4MMY2P\ZJH1_RIB@D9;^H,&APG@D>RT1dNg.RGgM30bKf.RSF+<<)@a>87
FcZ:=RUX8F+@8.JX>/d-eaZ+K<7SP[#LIKDM:TOJ^FW#GMX^S4\I]:.<93Q>8b?B
B//7.Z:;.R,0+YcQX,6]F0c_R2;NTbbIYIO-g@6f2#]B^dIH,FIfE6CPa3[G2ROf
@I04PYOQNB;_e:O8@e7>aYYM?Y,EFM+SE>/3bIUPJ/OM2J0PN)AcRaFZC-UcFY;U
Tf>NQPeVgGG@2c64>9ZX/cP^F47RRQR9aLgM&QP04.0?_7f#(?ZPg)/6aZVNCR\)
QaDZN;Q#e+:\),d8&[JCJF[\A#[LU0P&Cd1?/C@,0E+Bg;5<gb,)+gEe;MZQ(gNV
(2\9KL#,6H)Lg&+?_C<_/7Uc9(N<ZAOXAXJDF1:(LH.B9Q>)J^/TgY.+DI#I/<^:
eIH482ZU00T1/;ORROQVK^bAKVDPa5)=Me>b/JbF<AW@Adg_deJ&OG5f>OLaD^gP
RV6>&g1L:.<+;-9LWgc@H@9K4XH^UK3BL=O[:#;=NTQf9[S7YDG=(0,c+-J8B2Q^
:1\eM/f[c&-Me]eX#KS09XT:1ec>M5f&fV#JE.EE(B>KOJ,\?YB3TZcXT<^00H[O
FQZ^gAVdd)Q4PJ)OD)&,ZL1SQ3LY44.F8WNKBDbZNK?G=E[7@d-@G2HLaJZ>c:\S
O6bC1Q:Q;Yc:FVS_bb84a)RA-Rf>BBOA+,+1&MW-F/eMSJ]U&B=,K#;e2VPWK(A;
>^Z]6B?3ZDUg]QI(.+^A4f8;&,4WJDVG3/-#&U:fJ7\^1L7/GNT1T[PYc1d7C7_e
A#6SNQ7&Rb,FD?MD[A7f/4>],Ygg6BM0e^DO6@d]+/dVK<ZE)_+>GF#:JJ)HX(G1
>V^N9HXaODb#XPU_.)[P6ETg<dFg279DA[Q^.T7fd7/:/Eb5YR+b<dO&.9-)b+B<
+#.9TW2:\3VTOW&N>0G=&YO4AQXQ0Q/BHEQ0AE_Y_fcYT:2M6E=J>Ca&LUFgCVcC
I8Z<R>H<a//0.I-1]JZ\M>+VV05(;dFb4PFcV2+NT15^JBW>W#K1J:8eYC<Sg6<V
JgGNgPTBAg6RZ3V25ZKZ,?Zb]5JD_)IgD4Md.<R,E/D]N8@1Kd5a2,637W_9^2)T
Y.HDB\11,+cb\<VK;)f9a<>PFWK_Jb4gR>GIS+Q)VD<Z\&9;)#aEc=P94,Y1FKGR
K6S&E.XP0a[g\-gCIV86W:=,JRBTSG8(O5OR<9&4f-D)M_)c\I.RDK4bO3A.5N0c
B:2USIBHFC0FP)7A7RQR_LQa5@I/N(S?;FT7CVegA3)?GJAE8S2Ae+dfOR5AYbF?
ga\3PESOaFMAYVYa3X8R]YBHc33=,Z<24^C)c23Of=6G#Z-E)R52CdU/J]fb,S3Z
(4J6RU)S6#JXUPb^@dcf>g^Q-F\#>-,WR:e=.@Z92,[ZG&DVN<7AKZe/E0_N6HaC
O(:VIcC84,PDBPYQgCX,baM_b??CK7^(]4a+2?RB&#.-.Y76?&.N]?c7;U_CCDO#
=<A:#G9:gN9Ab.8?I-d:UdbGD4;.Na)\.GOS<7&O.abI@2b/9Q,23H>[J#EPK@C^
SYe7-.LRe;LMaI25Qe?b?KaQLOd\LHJef3VX\B=F6)EBB:[<V=9JY74)^3RHV[C&
gD[.c<E4F\.D2B=c7,>CX)RA6]/QNfD,TeXRG0/YNV[(4G=F_B7[M-7PgIgDd6\b
[IfX&5@d7@#(SU(ODe4<89(F^.B<KYZg8/?f<&/XD?0CN5AebJ>?WPB-(=\@CP/8
TBgVFc[-LR0LY3(0S4(3M6[-5Nf)62YeT,=&CBEPHG.L/-g/P/L[I(^Y&CAe1\X\
<Ge.N,]U9b#=L>gV-[#?X<d86aB&Me)RJS>;TX[-N96>0=YDOE+3M/-7COce-L3&
YV\T@b((F>21fHYIN+<JCg2;S5PF<<<g^YPI&Z4dU]6]9]b)@NP4Y[S14;N\Tc?4
5a6Y5_+(S-4W+<3_X^8+3gH_MAKRP6ccTGV_X\]ZYfgOgWR84+\.F@a15eGHAcUf
[_6F-T8>]@;fOI(LDZYNW2gfde8JDF1-9YWfV:2MP.&&Fee?^7T0^RRG,_]4,/F2
C354Lg&eD(Y,2.TU+]J@cA?,CV3(I9^]U^^76)8ed:Y]g/CA@\=\Of3JUEQbL8&B
E)]Z<3dV+E4aRR/NYRfN6IU2XF#8gMW1OD3:EYeZEN^XXbVQ_aT;^:P;MU2)_\c\
_XH72;IK[1@:N@IAM:\BPCL5BKC>=DV;]8bAda^)[1eNYVaLL[\cK?cICXL&I-]\
2<\?aP1B@6QAS,4[e35DK(_@81IDHK2#Xf3<Dd6fRJWa)+;dg+7AFCE<?HVRZ53F
8U@+T(3FJRcc87K,c8@?b\PEKD._S2)b^Te6_CYY1b?:/NE_8E8.U4G\Wcg,P/<X
]H&?XJgIbY><?N>WKQ2OfU[OULX#45G7>3FMXV;?4]TC-D(VK9X7C?ZZCb[0OLFP
CeJ+KdZG9<)MT@S4fSDb\5+T_PDT/[V_KD=-^NM@(PN<C1f=>F&Z51;Rfb_d+^MF
Sb3)C<4)5>Q3;ZFNdFQDP:<X+a&=ag,\]KH=4FC/]#+S]:8V5];&ace&/ZB?WFL\
aL3[PR5>=de)G_aT>dfWa^d(6JY^J+77.4MD4)^.VV@Z37P,Q4WPB:cQND:\PTe9
_DZKE+5[L?9?V^;L^dPMJLL\HdcIIC4cM2MF/dTMIEBC=M.(L_#KcN]CNQDJB.@[
1+H=<f4OAH9-<O=P72]C89;6=^M(,=,1;EX+6bB_#aW^fAd@Q\eA(V+@Qb72Vfad
>-,Y.E<)HO:T\-G6AP)GRRZ\LfI7N\5@M9F/ALQ<&eTWZPK_USN&6F4M\D(B3E5X
6]D:Sfb:X-O?=UNgZ)://84Z-PT8.8c_VUeXad^Q15<beWfAZK>5EgFF<C?5<7g&
0dK5<.#/:.&.eJAK(e+,,Q5#JE8QU_IV(3gVS85RI:e-,fZ&J4eMP:6@/PI0,1NY
G.Z,YLf=Q\?PYL6=_YEGBaZI>5X#AR-2=GDMFM[ZY0ZWGDWPWKf&[?0M_O#<>N2Y
5CbI>E(fMgC9Xf9]LRQH^46Q=M/a;N;P?aRd3><O4VJe4,BG=R];P+)LcIA8gBbT
.YG_)/Y;[\Y1PZ#8)QS,g#Q1>7?Q-e4:9#6:Ua@+RGg_UEO0\b8fYG2)CQ,G2^RY
4VZ]8f^;baaTP-\8?JgO5/Ef+e<8^\GP\:Ld)KWD&,(?U[(&WeQA^>d\W+0<T3(3
5C([P5<U(O#BG7b9PS\8XPPF6gg:ASL+CGC;bFKWf71YMWM&AV>^FfZ-XK:B.XR8
M^F<?,_e0#+H@C7:dAV9B\eN.J@.fZZ,eD9<C3H7][XFO3V+_65IOcMQdR?<dOfb
U-#24aKQXUU)JbHb[\-f1_X5??G.,N[X.A+7gY:bLcGO4A+<e2Q&OWMZ]CN[8K@^
f4M:&db,;I@+d5:f)XU)fMd<P)DP(KTPg&_LPd.B;Y7L4?0(<()]UZ?AggBQHWId
<=0d;LQ?WgJbH=aa0S:XgWSU2Y.F6,>R:??AN-9O85]Q]D][51<LJ9&PB:^NDXX6
2WPCQR)G2P,V_XQER<WP0^GUUN2+7eK/>F4>]7LGc>gT__0bc]=dH5MgX;6C_T.6
N;MU,RM7L?;_?9;?^-KSae7U_aRU9PUfN;H_7\aFY4N\1fM?@b3GI3eaI6-]Ygd)
C@K-36/2^-\O&JGCVI^<(Y>dK,QT#Pg_\C:2fVP=?G+2BLC4;931P#LYS+3S<P0]
M6I9C)]2L42dIM4]HR1WF[;F/b,8f1CQ6PYcE;:g#.,Z<RJ+&P8_D.-ZQeL(L:0@
Z#<X_2[6bK2PgSBD3H17)/J+676<S=4#(.E.>D(AeN;R)@69=S1aK5O#ANZ8@(KL
R+7G@>4.EgIZ6S+X_eO+bARYIMIS#W5B@01.?R]fPFR_1b9PE43EGfaP]-LME:a2
8;ZYDIeecKHdTUQ56XP:OV9HGc,(+NIEcbV:0]]OHQAIgE])3aSY4c.LAc=Z^5WE
a<N:6X1KVI]TRT\D0M^=a+VC50DK)+J3,8d:M3<]S1fPC2VT3LIH^S1X>QM(>])P
PgY7[(4QP1CDg>UYJ)_M\K,<W^aS;?I+:AZ8NcEc>7]P..L9,^=RfX^DP)<O#J8D
_JRS@(X_c#T/CE.c\W7W0IO<CeU=D4F8N<0,S()3Y59;=U1D1H#-.;HYfcME6Q-L
SBCF5SQ99ZJ_5<g5:.;D\WC0,E(J-1&)KW,&:eaWRBP:W5E4^a&c7H/4D6Y;N.3_
;#Eab;IDXP&RB<GO,gZ<UE;=6:#aFeZ2.0X@QN/eGLS=#>UN;aSc:<GK(-,Va[\L
=4RTb^5CGca_=M9:>Y.ZVQd@1TOT_/[VcXR@[&P)^_HWLd(B&5F9-)?>3<=T=a<=
Xb=)bTH@<CM41HG6O_eQa4RDf<<_COO?<IV[]f4IWPXP5N]H3Jc(_ec:(U=VRg4d
>[(2CO<#H;\#D7M-/9&]Je4TDJ#V+KSa@09f4G&GI3W]M0Zg;ad3:GQ\S7N.YZ6+
D0;8?5@^;,@XB8I-#c0#d4S=10RK84e4>Aa4-_3K9_36Yg12)=e11[T>H@BW;X7M
)#d81:EPL6IPC<^Ue([O=MHK]S.V[[bF>5RCME<H;e8C0<Bb_60d^.S\,7cZVabZ
WdU:HR=9K>V?\dXBG[6).3;-46.^07+W=^6FaV;)e]#]gd/JdO=PG-2=Mf47&(Fe
79EL7VZb#[G7/DX>Aa[X2a0A268(+U,V=ONTE)@6@(Mc2XC-)1+>C5GC68A_-8^E
CUTbG+@8XTD+3d7Q09-eAL.-:C(]53JOcG)+E[.C64T7:Q/6VQX?YKV3FHBS3;:M
dBCQD2fEY5)<T3bOOPIN,\C]0VX3T++<@(ReLP];a9C^@HR/77>A>?P.]=88+^Qb
b7S\Ef=9;T:L>,>_J,D.O[7a82&#c->TUKX7eEVZ<3=1[Oc?.d]6X2F9/T[fO6OL
(KMM-<cCV5?:^8&WU+c)>B=<F&]))B1L+:,dc(VU[JYDC@C>@fI?0AU#BQ?LD)?8
U2^0N4^QXZAF=+EC#?0DJ<)d^b6B79U8=U.IWJ5;D+ZU[\.Cd;U/]Nff<J74(<@@
.EX?cU<agK:,aGa[N&A:D3?.c0L;.P5X.;S8CIEFVID3;a)87P\@P58,I\eSbDI/
C)_.A\4e@a0EbOd<.=-f@4aB[37,cH.&R^C(dc1]G5G\.F79?YP>9eQ3@96:()8g
<g&3c#0b\?RTePJDbUAG>5>IQ(.(9e<VSC(7D[M-+^YG4aYR&e<9G^C^=1E;.755
-U9\=.e<V2B=Z)<9dZJeC9:0<>>XACeTUf/6)6/Oe3,;_e.<AY;1O,Z<D@+?G;C0
f:M?6.PM.Y_AJ\W&S+UX(]+15^b77<FPLMGfagE2((>ZK>^I)[9S)G6KDGE4YU2:
g22aA:e7c#<\e9E9-QWW^O]@BO8PF;B0<Cc701R+6M_JG<EWL]R/7W7V>P/S<GLC
7GF<U3=A?gP[;KQf4Q,e(,JeFZG./gH>NCK^IZUD2KJ,gD3B6?2CQe0,;BFcF2\3
WI\?.A(>=9L&N.g2_g.D3I<.N/e9,H-?_0-&:LSBNZOZ8V@9BR<I:K]UQUXD5::C
bU7PI81Z\cNJ/:H?D\1:7H+,^005M1/3^JXZ8RG^B:eKJg)H0ZFFS7V)1\:g6d#@
P.4Y#VMd40_4+aRI0N[(H0d-MfXLNd8fX+P79KF&XbKD5O,PSQYIbaUBLM1VP6@f
b-R.JbDZN24]S<T.HYP2(d+f]^0LJdYe@#R_CRV]Z+PX&K0K&KP)gGGFaG.YN[6C
Nca1B85?>72&2?X_I]GX).RENOYe9P7J)MeWSHEZ>_^_)IRfT@/N8K3P<K7d0bNP
eZ_6ZR(<[(d[1,UP.W.eQ4-5<IC<O4,9(]#.MI#;BP>;;6H1Q+LU^6O^:QVGR1H1
KAA)N[B6EA7>BUY6&;R/Gd.1GBEO/:=@^RFNU#Vd1eeT&F3&[I97GUTV+XPQ\aXP
K14/-W@3Q:T7_9^GfE2FE8;W5()SN)CD(DKbR27/KW]\(F&G.Sa@B^]VZ7Z+B,>;
ZR[G^d[EeR[5CUNM6;Q/ZEd;\6XQ@-(gQR,__@c1SZZO\Q&\c(<Q-U45GD.N9H+U
.JDB38CJS1:V4cCT-V=Cd>Gf3MQQ=B17@W,3+M+@^X060:#:NR/U1\?=<P.>Ab.=
f<PTJ+ZG#DS12C>-R(E^(I6Y)+><KQ-A.74)ZJI/;(>G#DDW##QVGeXI./d?2/AM
0(B\d6d85\U@C6;/O4/=M??aWU=0X9AT433HffBGUM0(0\6F<Q[4KFCdbf2^9>/.
R)c&UD,efO4d@,:TZTR_SSWP[YRZfWPQJRYB(5bU(&Eb.>MDaagKPg^:@P?CUZ(d
\>;A8d+-+,=T7\]&QKM^:)4b+J9e2BX:=EPT6+cg@=&OTc2I.:Q)((eE1&f=35#(
#)I9]C(BaNYLWgUL:T,<3M.[Mff.W1I8-5G?0O4c3?OM=)PeT9>8\O.Wec2F6a@d
U5.[TAK&0CRXeZDB-/TTI[NRg?JDLFIU:0OJ3+OUM.b7XQOQ08<HJbQN\5dKg=?D
H.-MU;K+B<]=#TVOd;cb&=>,W=:SPRLVXDHJ_8]geYQIK0RR3e(A[>GY1=EHd#Q7
5/UGSfgM^S?U80J/MXFRFKJT0Z3JJ88f0CaIP?Rb\2K(.8f:YG#H=OC0_@H/;D1<
L96OGQ[;U4/gF\D0c(1K#5da1eP?-?d/N0TN2CU>K:)X\2;>XW4AZ>[>g\HZU7)R
MM\Wf#d]FFNE)W=8DaN@W?E)YQ@Qa#;1L,V^+NGNg\Q?II7&3>dg=^.[NO&)Y6F&
SZ3>&?V->d.]>6G+)c]0#,,fN4NXHBWW7d4?LR9Na/Ab=5:BCfDU.>P/FT+6>-)\
KFPI7NI\ASWFX15FW52)4(U0IfACK./]=X)/A11(8VT,Y#R7=OA^P?6^0Q9HE(Z)
]>;BLZOH24(SIW,Y(@?YZHfHJ_7W+dcX4aGJO2F[a?PT8QY8.TZ]_:&N_J13I)N3
YV7a+>DfMeM73J?G6CB4a5FCZ9Z4/aZ#O>U:U\:b7[#]5cUY1F<TQe7D1bTaDV2H
c\<3L-.ZJJCaGFCI1&ODP6Q(Y0FO+Zf?;21\F)]WWC,SNP:@X^WL5-/dH@eUGX)d
?QLPC^65?PWO>8^5=)<CRP/CR/1gN5I(OAQSMZ)>2gD:O7-G-;YbfeH^ZUD1D,^&
(>DR-2T=]b1RN6(bYBAC(7\AZ?J/NeZ80RNZb\.[>cR@_9)&-b-&Y?GFbD5.SMZD
O:4J[R[[Q]fF^CgCMW4T]8ZFAY;PcUU#BD9=J8M<9a@);H6d<#Va5B1<.A;33ePG
?+OFf)4^[(:W2Gd?]BDC<a].ZBIXR:[=/17BSQ;3O1ND3YKBZgF1)4?,BJO94MIM
Q<7JYH\0E(,U(f&I\LUaZCS&,JLcTdc]Se9<BYEbOIJ)X.9?C+.M(#V,M@eQdLY7
e2B;H(C>cGJXE5BO?<#QNT@TZ,)T73Qb5d]DB&&Q.&PIQ@0F0XVQ[+EQ[=)BR<UA
eAfK>=SM+a:-/OB5UJ(B([6-&WF6D[ES?c@d#,]I_4&J[KH&_;OQWac[3dZ3c&NH
)W/HZQ.MPZVA.8H(NZ-d_E/AW071>eINT-REY]TFaZ9A]D/<ONR@V7+P6QR_P,YT
(ELN<S2@V[e94#0<&^PG<.&AE7c>fM6>I3B_R3,UCJ[5F9<]LS)f1GJS=G@O@@)R
:CCG:HV[J^Q-.dG9+8&dZS3M9A?Vc8K?IaQ1FJ,6d5YHY#g:=,dH)7a2eS&_0UF-
e)FXD[.JKb\Y(:VP\L<-CG:\@^VG/R[J9;@O_.UMA0<gVb6AP4;VH+LDEGT9^[-U
)W?_]>5Z3SV+#HddU[^?X/K)@^:[RU?Pf34K-&5g=f4g[H#GM\?XZ:8-R9aYGDM)
X;dgL4:40CdK@#F?:>51;e--;XG3B26-3dBcSQb#:bWOP?+AIJ\^b0;&[J=M2NeJ
X[(J9fgS9adFOe?2f.9g);)B;-b9f#@N0S,&GgG@Id@\-bgB(?b9?g#c[)ELc(eU
0D]J.CY_=3UNUR:73(VP7O.H,#+3O3:f^RdCFVcQT@E]&0f>/DG6,X#U7#/=7.3a
7AR&@UWMdD9YCW]\B_?W3@CFe?9B8W1?+BZCSAS41].VdW7Je=JfTFO4#gTQ(G=9
<f:])57>)?+7#cd2P.ZQR^Z=GUD:Bdd)2(Y<^=MZ3,gc&8350.9gY@bNN9V,>e8Q
=5V3Wg]<KE/>:>H<T\>6bfHFgbfaIHJ_EHO0,001BPFPXCNK7NT;LO_:QRJ^1G,)
2F2EV4B+Z/I@VdW^D?,FU3<WfFRR>673FGC(=9)IK^U>4OaZX(3eCZfP3<)cYWca
(KQP1\<-I&;]Vc,/:+N+&bE\QPaX=d-^9f=J]4=CD@HK@P#WQU7bdDQa-&@456B0
5C1N#)&?.GfMZG85Maa._LQf5CRFI.J)?1K3GO\/T1ZRMX48.J;#?+N/L:bbJ/0_
+@/49RH3dQKCVX[aRY6;bR8Z?aQJBc^4_Z?B014R]Q>^\;(9N)ef#6Y=RdB\)Sce
DgWLdXSD0(W0gA?8;&6b9M-)F8F1NZ5W@d+b,^+PG@R#3NQ<13?H+JOcT5Ef.0e<
HSDP@V-<W)WW_,d_+DT/6GY5b4J(3BTX=KRH>=b]O2Q2GBS]KcJZ@O[=PSZa>G<a
A]4\-/BY,a+Z]^.dg&f(eJ7O4\N4GN:Cf[--^(0g[ISNDg[b+,,QWVJT_/SgY@C?
RQ+X2^NZ;)=D98/]/R##]CVbJ7OJDceJOZbKf9Y;e8MbgM;EXWTFWFbPASM3+&3c
\e^MJ.GQ>H^+I#W/-W=)ED_UU<CDPE;=4IUOX9:C=S<(ObMaOaY9()#9A,RKHW(g
Q?.&>gEE]U&56<)+\K)+P3KX#73f[+?J^>0P-8TIH:d4K^EE39R]O1JRR\@A3.C/
9_I5#0&fZ=4D?RD=R0\++O,,8Y=AaFXbLY5O>?(D#+Kf/(SZ<@,8Rga,VJE+706T
e1=c<XN[>T_+DOJF<8)<I+T)eK+5IT;gC4,fd^J&(R.PQ-5J<UW9Nd]D)@)R:[;(
?Da,XgDPa6g[5\g5V^KNT6eC,R99;Q7W]KUXDc/H\R#E4Vb#KT&--/].N/)H7c)I
_HOV6[Cg1Q<G<]>dXa=QA^62#LRU9XK./\,V5/O6)5f0E\KJ=_/38HIUKdI:db<b
MRg^?J+)E&[c5GQ[4NF((#3:XXNGW\Jg9-Qf;IT/R.J[dbI\g<^B6F8-THQLSPT=
,a)-I+:I#]aC/ed=RNX\#+CDN,0KH/3\YJJA20RBPce-2DCVIG8>47-O7]8]dH4C
-H\4dTIcPIV8gN2P.VR\3_#-5dKHST^88a?74bKLPFaB]GR&CB+a+(gQS1-OD[&d
aD,&SE3(da,Z#.</AD(1T==3<\4.V]FV[cgVM]SU\61e-HDdEe<T/H,cH4Z83)VT
[HX=#(N./=719+6K-;c)(7/2.[,K(A&;bRSDeXZ:1eCf0gI^X,BYaDY9F7B4M?ab
;HJ[>#&SQcHKVH7]]bH@Y)4)NL/a8_OMbM,99<EfG=MW+8AG,N0KQZ[<LW+&Q3:;
X[SU=8(fKVgN9A_O1(F9\cLLVbF\)RF_N.)ELPY=c+8+HZ.dbcSaK?P:MVLCJTDU
IZIEOCDGA?>9LJ#C9@JN\A3;IH,S08?J85d\9C?^MFEdD_d;Y,QT_H:(GJTabg#J
GeSA]RYfbCgRE)E5<;2]5a\c1b:UF)BcP#O,+4Y-E2?L^>0L#1D1<R)af:]XMALX
<g+[S,\Q^,dHGd+S@CJB49E4c)A6FRgJe:7D&Z7&AIV)N4.X5],(4LH32Z#H3A7f
1g26J_BaY?Z<8fgE-)J:Q4<T8c^+7V^GQ9X.EU)>c06(UFWU=JZ0Eg+\c0I)^SV[
KF9876f3.LTg[X=HA<9ZGU5;_@4>3QCV2L?eHg5E\WW5e;8:3(aL.&@/;,@I+B;E
1fSLfG/(g-(P+-&Y&-PRQ_T<STfY).71U=M.a.Q+^/ebJ5GCD1Ka^5=c;P#[-LZU
+IQ=0?/>F.]BON\A?fJE>_,32FE(6fR.c;D<U/[+5[8HddEHF;9Y;RWg:FF\<R4Z
^PS8FN923Zf3A7__CG_I^LFR,[TT<eF>+@7,Z<[GgKA>4(W@VYEDJ<5LP#12=?.,
=)/d=1M4.I4cRR46C50=.;ZGc9e4-M#+02E[^.(M5L11dF2T.=6NZSML<40NL2L;
=-F]7@D9aND?&b0S]?4]8\1.2d&EJQQUSD#/0)=[_332F6SU?CKP5+bV_<H_50-Z
L;WX=_T,\S4U7:/YPUO6TX/[,OG2YS<-U[3a\b(3>cU>AN)#JP25.79?#/1;bgL-
?DWa\N^/W]OFT3N)0.Md7?>LSFebJa_)4;WdP@/8aU@+OWg;ZE8Ke>f]bG4.L>0?
.SFa2(P@a)7IXZBYg<?fF6PJ9^ADV)=)E.@d3Z4[/4fEVY/5F2D5(DL?>7Ub(XbL
,:CHfTd@K5+3+@g?H?#1ZcPN4-WS&X.Z=0RZ^W\VDCYW0]TO_U(F6I.[I>)B[+0:
e0J?I@f,^:AZRF>#@Rcb1,B^0RCgAQfX2_N+b3D6Y\R2CFK/FYUQNJEVf[87,Pc3
e^c&:dV\,PM\(9M>&LQ08))@L\G/1,60XL)4FZ:V1PKf)dUbFabD2geC7AK030+_
?<J75aMe\/P1LYcaK.++N-0f2DF--=f>b#&d@Yab^V]<R_8/YYDMP4QbbKEFT?RB
](1[:I0?Se?]45Y&.MI/>_K[]:RW:J/@K;Ye8IaAQFg##d,cEeC2:\OEO]7:b-NJ
F:.-^0IZ2X4f;\D9ACEHCHaE-WBI>G[FNFZFNQFDgK?ZJ-@>URSLbXWd@G55OScP
5NSLVV3KB@(^5TY^CYaARX.=N3>HZC@C(GO4a(QJ&4((0V.\4Q:_15Y1eSC?E[=2
WS78f0@W;HWR&?<8gFf,0POb]6TZQ5^E5^X.fdI=227G62UOIG8-#(F<KaIVAOG#
c8B_5;;,AWNQ\2^]e+K[.FRWA1aFA(92Q47TQ65G27HA;O0d3/fPJUPVO)We@-HM
[17BK?PG^YVBY)VLe4PKYASTI;^QS^RYbTDDMc6O^5c5-O8R=LI7:X@2]bRNZOVZ
=feL+85Y@J4_68YCM>BKA6XI.7F0U4;g)0LE)e>a9-/7ZO]H74fe-[KV-_Ca/5Kg
N>^22ADW-H@=PBO5\,M,(7?SFMW#=-NC7/T;O>CPLdSJ-?G&+a#K:Eg.ER<RS/9d
-C675MI(J::d2FH4Y#,P(J\X@9?M2<X/:[[K<eSB+Q#QJD^<7=8cH.;9:-?REP//
XDZ0<05R&6=S<-24gUMNgSAON?FDIL[]7JI,BQJ/A&+P3/\\A]_V)ZbY(:UR\3\,
_g&[=T29AG+=YM-RSdVC)VcU>0a_IM.HgSVFV5cF?^O0UffILLfRd=aAVP<HNZ-6
E.7P6EGWU?H6eFb#g8gKc5-4.=3#@-38#+c=J=95;5]62K4d,X7UWL8>#CZfS8G;
X2>2>MVHC7LZQZA3-(;5[V00Y9bPd:Z@YKNSYff#7[A_N=BE0=g?.4S#OT,0QMgb
1A3Md1NM/(SGLK[1FE8&H3HeQ=cRD3<AQ+F+(F]YdY0M-&#8O0#ELP1:<W9W]V22
>cIIg.d+R3Q3f?O#I\ZJF)bIE+/0HRO5T\@L.7@cHR?UaWADb(5<HMKY+ZXRS:JW
=,]B7W,>>@96S&(V9CM:L_Q?a9C>ga1P9IM.II-+1@:b_N=^5PLIE]JGSWT/)FLS
>Ma,7Rbb@HYXaO;79,Ig/dKe)S,QLK8T#&)T5]ZYe^GI3E3VKJ?1GD-GZ,Pd?_]C
@?7B=WBS5K3+g]<[dV:2GTB=</2@D9[4;J,>8<R8\fb=/7Q4]1U./+bU0(5^KVEB
3#@g;DA_aS\S\,YD.:+VSd8D9F34eCC;:+SWQ-TWYFPI/NJ#</gB3>J0:_]VOP:T
.QD5OB@b-IZA3W+(86fTT92L08[&Hc)]=L;(3LZC3b#.__LI-8C=_#d6IVWEQ@V5
FB)4)dST&FB?;;X4X&JJ9V@c5fV)1R3\B4=1=QNESOXG2E^dW-H<<:=7e1/O;KCY
/YL;I6O=6)F;2HI=)Bb;Gb1bFM9AWP@O)\.3R:GP^[e/D&aH)OK_]D.HFY)(P=E#
/^O+WEUHZdMN2d<XF7\TP]2XQT2[BJ/^;@U9gCZ2KgT<C+3eDdZXZ.==UccF,J[B
E7S;_,7#bTC>;4KZTLGbTP@>G>,3bLF968#D0fVE\P70GaB98dY31#+(46HDQ1#F
7,gN6C+gfH2O?2aU;:/??Q=SFe52L@FfQ3_PF.G[(]43<C#ga5\:18U0HFGRXb\.
PS>_7.(00J2CMYQUB\,b-<b+<LO)WTe/&M[8-QM\b7-J_8c=.X<=7>>I:YC9:d5F
7Xe;2+\5F;L)@1:XFD<O?^Q)FEKW9.a>Mg[-H[TJA.DbDLFVJT9f>F>=PCM=^=7#
fU5A_L>EPS&Q2\aFUJ9\&F#[a21UDW@5:7#S+bRGG5:PF.XR-G^RJ9K(H5Dg\VGU
Y-;>(Ve.?G&52WgL(84W=N:8_I,>;=K/g+K(<D6aOH3FQ@a1,R]-<SV(@8X;V0Pd
OCJLfQ_(^_@]HC6faU)QX#VUJQg-EgFDX1OCEN2_#VL).2TJ9g-dMY8PU(>25C2F
YMed/_DNDY)]?[#@.QIJT1P(;NTE4>5_fbYcL4-fU2PfB/8@+_FBFJ:1W8AaAKR&
#5Y]A^d3IYM5DXHM9LY.)0de)(IE:PE_UP:T+^B.7Ud\c;/P<T[f+aJ=2VF2TV[P
L-2<YU@g:aR,CE]bS>=PL&BgL1&dMYN_F&U@,34R^?4?eaeZb<Z.9bb#>ZLbWf:N
+KH9cdGW-cWg.CSDTaZEgSbX.<ZASdHNZNb@7P,UG33_E.3FUf#_\-CE]LOD00DM
X&B=D[bD0OOQe82EN(RIe<=O6C+Mb2Tf(YO]fU^GGEY+KcB8@=XZ\B=76RTT=K-P
_NFP14J]2+BV86:OYdXf-ZO==F:FfbE-,gBWRD?TOeAP;Z2:b/\94U/53X3)Ub+V
)]7\XX/bCMJN1<D:,3K[=&+K#1I/@,SYU)N7ge^]?(fa[G[ZD\IZ8dH?FJ_/P(1-
Hb-_=P>a4=e(8gaCD[AXP+e5:5BL7/@#@2]=XB1DQ-b_<#P[[QNC>(2W&HOL74dP
Z(0-8dO<\7<2>H55Y=8V.U<0bRUZT@Y&2&52e/dF_ZK-&g+)beB#(0[c@_KF>G?2
:\.4-cKQ\E<H^:-2;CLDQ.Rce;6G1g]g+DE6?=F):E-@)Y;Idb)GL3&)d040b^^G
BXVFB[g1GQ0c92),CW9I/5XG;,]\c5/]]BC67R>O>Na06G1W<))APg:(40N-/^\N
PEPXKR0?A,ea_aI^@A+14J8L6=\C[,1_4SO7:P_/R>PQC(UIcY(7OZ;(U/H,42cY
CYZ5TNK7U&:^JbUe_a:e:1X8NbR?DJ0ZXU4b/0Y;b0NYLVP]fA2V@KD1&[W?cN8A
T]WX;9-HO.H60SZ^ETYY3;;I=5VT_<0_:^B\;)f_eSNABE_H/X0AeIXe8QR8C/+J
2E,9-BL&:PVDOde@OKCeY4_fHOgb,TJHGKL\GNZNHU]e;e8<HMeC^474(3^5NJ[/
c-K<_&fNCC?T;10ecV3_C9RcB_3,cK>_[\U^5K64=97I;Zb46&P5a182A699c;MV
ZG&MPV5c#:J0fbeT7F8e^;JVRQH]B@@NPMTbdgKdJ=\:TK>#O0HcM3Y432(DHb:\
SA]/S<=e.-V=3@(_]Z<EI?Q&WBND-fJ>e-Q>W=)8MI:LMU&cXC@1_7>HP^702P]f
Ng2?f1IGAP\a<e:O/9>2UKFHXXPc:5>/V8EOF4cXTd.^C>5GE9+\aB5XEH]>8=?8
F.Q>F#=,-O8NL3]81AC@0@U/aScX+,JHL5E#GafD^V+B?@a[65/[67aB;>HX&ZfQ
d2#P4O3Qd+(SeQZ\g.@MHZ3fTZfSV:aXBbE,9cK3A7VT-d)D]BTIfbNPIB_OW.gX
&)Q^I7@6Oe4,W79-CB;\/?IK7Y#[JL+S(f0SD>a20XXYP&KL-2Y\?0fd3BOf8^4e
<:W]a:MZ7a8B)&9?0F@NAIRH,J3^c@N=Sg27@6X;D#c1]O-e1dR@.A2>_fd6;I)A
B>XN+359OY?ZJ&TJa[IR5R.P@XU=)+FbgKc0?dJgY6gVVG:OW^]0JT\;-(RC0aM)
ab_(AJ3A?,+FJ-&8OgT05cge;/7<C6aX7/BfE01S,c_80;3/;H9^4[Yec,-5/F>.
EIJ1?59(2EC8^VebR9M&L(_(7EUM0;SCgFe;fJU;6M;.VH-EWS_T8)CRV/_1V8J8
BK^3-&UT382>ffLSe?A+\?ZZ>89[Q]d)X-=--=7]IN@CA5^6<@:S&6&4IQ:KK8NI
YS@,03QcG)7VK8e=EAG4R(cD/0(+fQe;1NM2H8_f0S.:7Hc&b=T+eY^=(SGNEO?2
B]T<a./+?P^.0VW5?;a\NgB-@R?;008S9W._RBJdbCB2IRga6K._6E74aR@969^g
D3>BUD5V<6\#UaBHOH3beRFI=SX?c>dG58RXE=Q3FZdYZ](ZKAP<8NFgNX41WC/7
+8Q1;5^2Ag+EGf:(K[GB07]##-5dK:;O9(.DN[_:1]]6C(NRTJ:I8M\P3P>gISZa
W(SeW&-[RM;g;fW+W+0X3TT23-HeABfKPR&LK:YV2^()8d,@411@+_-,GDVb2#_7
0>>8@A5+g^[H&ZZ(XO>1c<_g>LOYK.EEGg0@=.TI+F-(\:6<a?P#_\0+V^a^]b+\
T-R(L99;6?O7KUL^,b_@Gd@)C]1ET5/4U@XTK?G<3\GHBL2SEJL3J^]^U=\=2Teb
f-LEc^V1D&(KggVS;SKCE_O;;EMBC[QRIP_EM4;RFM_=Ve9RY[7+X)3#].(,bKF)
(1D6<UM8aaB7W[\J85AMQbTXWK-U>VEU]eAT5+TGN1dF\7<]O\MReW/:-aER3aH[
N,,VD_Zd::N0.PQB7Qe5;<9[6R^.7d@OJfJ1&(VE016ggb,g/A;(E@N@P)=TG3NN
?IK]3X3GMR_2C89JgT3<f\K(KEe:691#;>.MRPCNPRHP/[g#DNA37VI6e5T/<dW9
]D&63N/Q(Z)-bdP]L62ZMW\@BY#(VG^U?fff0gVbP5#a\[>TA9Z6H6X^5>^-I7@0
.G-&I</OD4,<3@>:HR-P_):H7HHb[#&JCHJ]HDcUb(=:<X39^L+,>(&-7A5]:,_?
VKg#5OAeF4=3?gFW7Wd41RB-0cEZTD9Y^UA,42Sa>aSOIIQ\F0L=I.[X3LZOOHX_
@)g&YOX=XCaX+7/.?3aZ_=NOb9Q2TD#8A@^+eO<:AeF-RPD#c/CEM8&UG3_&Z(_d
?><PdTV,R=HXBUS3cYDbNI<=&:A3#d9@D^+/g71E-aaL,;Nbf]YM_V51aaG#XHD[
/,f/4C/JF,T@O_=aN<eJ4X53632gIO6<R)V4(84A6N]H^4KKKQOO&AgW+ddW>+Bg
Y1:^9cH/C=)467aL^TDD/XHG#-724401KLQAg-D#,J.c=UTO.K+=RHVPe;=a1U,)
Y_WK6We,Y2^=I^D,(RJE9<&]68]TX;>-7+84Ce]YL6V5gG,X]ZUXL6V=caAV&H<R
H@B.Z-P3PTUI/TJe5MGbfT44R9FA1Z0#&:5F1,-8T,5d6H(^T21e/=H<+Z@OC\H6
-PZ/^ffPg1B@MbOZ2O)gg@ZST6-]QT_X62#9g+<\M\ZZ<S6UX,\MI6&\2T2L@B#Z
dSVSW/IT,_GYG<JUTI;6Y91);5;=:[gME)gDLKOQR6\9A/38VKgDJ>\9G:4[0H[H
\,+97Z-C;NEB94IC#@g=:Y=UU4<cF,PcHVa53^V6WAI5(1CgbOfK5MV>.S)LCP,4
:=X-f-]/Rb\UVb+a,B=Df04DRE4G_DH4eISJXW.C,<[PO9P<^+^ISKU,PL/@R<7E
aNWCYV\2CTX]8>0cCEGCEPC#S=>\Od+R/KP+(Y;(XR/10PH-HeA\0eX5N:c&I.J&
FYX)H2adDGabg#&F,=0#EDIDB?a;PeL&D-=-PPYeIJ?WSJUc5\-NZ4f54_@acgH]
2X+X_0JK:.@RB/HIA](;\DK)K<gH?fB/WXM2)._P.<A#03D@8CEfb#-,GCZYW2D[
C6LP@a1-&W=6N:8,>d4D7RGWC25+V+bI7)]dXBL>DE;C)-X86C8edM7HIDe#5=2V
3HMBCC;gR.4]Y\<a:V;.fQbb#(B/XcgJ=@^BAN\(5e@:,X=H02b,8<[f7#dG^5bP
,I#&Y&5S@PY3=CK\TOM<ab<B=Q?Ge1XU,P:Q>?9=8H+P8.KT@&dQ&aGQ>:/V)IH5
FW.YFKSe1AcJW(Pa,[)BE)NfN+f&\;@aC)Y7Qc-NWO9.6RX>ANZHBQ,J8AF:Ia&^
7O_>Q3=SQ-DD-JFPTJOBX8:@#XTfN/1)aM8A0+/K6(5CX\IYBM_^9/V;aE^W<db+
\48>-6T@A2X2>;H6WR0K7>NEX=F8DG&MQ@&3FF);_8=XWR/AL2Wc);7L6Q(#KDH@
U6INP[?b\/R[BS-7\(<SaM;6P6^Z;fcWSSVY].8Q:fN4I2bGa=)U?NA&Q4JG0<QY
@;0X4GJXa<FQeV[c7[MId-ZI1XPH/:T:LU08.EPaG-)O(5e]<M=g4GG2U/+[1WMe
<_>gP);?/7@^?:Q2IL@@7IeBJg,[R\UD;:>aVGHHba<#D1d:55+Paee\>PA/f#;b
B?aK10N#RI<1..LO:]AY)HVIJ/0.c3&#)I+KDGQ],PG,CX4b5:XOAWdB,<V-090]
)K2C9(-9&YZge[Y6<-JfSQ^&Q\3I,Y#1JTfNX-Q42R2_c)T+;,JdJ-@Ebd>TY/g]
X,\X64<PBCFJ153Z0;_ZCDMD^^9Se_L]WTQPX]6=a-17N:Vb,;8W4K)-cXSF7THJ
#L3e^SLXNP<E^fEZOE-FD,7KIOZ-\8UF@<GgMFf)Hc^0+fS\59_8YBGc:1D+Y4+>
(&9cBPFK4T;E(::Ib=d6S2f>;,W0;6R&<H+SaT\c+<c#AS_.^g]FFY;Z\>E9==;T
B:,9FE,]7C-TX]W]=-UCfV+C/JJ4g\88LG=>M3@aQeCXc2D:5EP_Qcb6[5]]BU:e
Sd=L=]Ub4@ZM?#D8UNYb;0Sf(:dE,8BC8dG@26W^##0PA4\&KV0K5GdMKS..ce=b
Q2RY)7AVKH5WMY.8(51<)09dRZ2De)LNId-L;G9W(VD)AON#BN@#1A&;]2?NS@9K
PO-.g6cZ=0S4&>2\57bT-UBVK#QRI8OEK0:94NY-LfPJ@ad8E#<9^1@Yde(K4OCX
W?_0ZDFgD,RfMVeIKJ.I?WeKM7@Ac>9KCg(QV\Fb?+;=;(.]2OVV?FP@+9Y;]Y;d
,]]FB2)0:822X=&2AT86#1)A[Z/E_SRV\;QJ<X-LSJM=@K664c.T51OVQ=2eP^fY
Rf^-?=Vf:(^4,e/S0a)2.cRdgD.F=EENPMZ9bLE+7IF]2T=c7.HQ2(#La6\3#I66
&N\0Wd=XL3.V9cB]>HN+V(fXUL-eCU=REC:7:cKHGK+#4[&]/X&=/<)IP&>ZPFO_
Z(+5:UMFb^]7SQTR-5),5d..4##QQ43,G+[YdM,MZI7+E)e34CXGZN#E-Obf2Vc5
8X(0JR]V:f,cF9_^KWOIg=f3+=9I1HX#EAQ9H]VD6FWFC\1;JU;@cR,c3ZJDY<aN
0PUZJ@^+=WW,Y^AO?TSNF8WQ=?]<b8X[.IP>3;(43M((7g1K=0eIdV,(gO<R12,C
LdBNAd/eCILEe\QO.@3;R1d_PHFLI\\0B[,eAT^5EA4?(B>DKVPW(9QP(^,<a-T[
02MEE6\8N/^cS1A^MPc-;g33b)U(A1HW\A2SXU;5/CMa6?S^4+YR+&6=]J=65)X)
V9.+Xg#/Y?.\&#STOaL]B-_J@;G4A<ASgX;Xg5f,e^gFDfF(QLIZJF^ba&2GNWW#
d+cf191\bKFZ+W02B^UBMfH[FQT-(,)<?F>_F/ZEAg^fB,\1^VDJ]2gf/b64X?c^
Y0&SaffM7=Sf@QD-4R?Ye/c2NCXJ+,4gR=,,P0cYB)-345S#1cPKQILcHXR4A>N,
OC/CgK,FBSY0a7gBZIAHSAA?e2KVV+aD+7/QYPHgFRg40fafFBOOE/D5[S+L->SR
+A3HJR6+N\&(-;7@M1G@aP4:W#U>LM\GKVfOBbQ0FHMCe&+c4X)::XFZ<S.E&MR]
UK9>7fa\ME:W\WAM?U:I3UP9:<Z]H&b\D>@WIFRXX4X[Eb0]DI@VeM:LIH6bSUI-
a4b5EL#+OLb:=TS7V[#K8@DT)(&A_&C)WT^\Jf21JZGUB;L#P)FO.\dVJW-AF.]D
WP.=P<e\-.C(MTaDA2a];b2,(0,2?O,>&4]ALJ:J\M/CP<XYU:faH.=:(Y1T0@f7
J#MQ3IG];J;QbcL\c?TIfXgN]BIUA2,;,Bc7U<6ZYG_2#D.9DaJF@RPXf>BO&ZK-
/F(OPZVbJI):P7SA@-F??8&>I9+SQ]Vb-65_V(UH>5WP)eH)e)(,XDR4[#.WMM#c
&Q+=eM#2,:FVZRa;/_MaJW/WU5C-UURC-7,f&4/d07ef\LOdP:Q5gZD]=;/+3:@E
cVY-;H:#PUcbLRCIN&HP8=DN0^&0J^g;7E&1f0,d9EKXO\9KAQe6M8Ob1PECZ/eE
/IBUJFb#65Z7Y;[K@\M0IYZPH=[F3bD7G>RgFB4A1JY\33U^G-JaO=]a=[b>W>_J
eZYc==A\1>_5OG^1PE65c^^R(/\^K<.cfYWBgV##Q-=e0;D23CPd[6>V+.?<C6,S
:e1<a8e/B\0D)/47DOeHa>+c3\b:SF44./]CT99XL03H:P?+Y;fBZFXVXAYFe[WY
gd-]]L33X_>[]&>U@N+3dX>LJSTb@Q-#CG_FYXEUD4L-(E_G]RS5_2#(#+6H&;[4
449KS-487.F,(aD8.V-AA)8(Q]HCS)V5L(VP.UZ71E::7SG9_XL4\IXY_5Vf)<T4
0D&Ad<Ig>b_9AF.,#308[#S?[a)c[M4F>HFN_4a4M?3-VV8\JN[;[-HYIe+.+U&P
\_C3XO[?A1A#@X=)#4V[-_K]NB0ZL@OY5I<ba<Gb,cW/,+_gEe[MUdc/A3ZJaO-W
HR+UI/B/4TW]BHUQU/T=YJHOX>g5O8R7@.[A6O\^I3ZPBJ\YO[N1?R&[)=TK8MCH
)1.ZL\f^IWX4ga1\MX_0/W>71YXV5J]I?,RMBDUYI:25b=D[PQ9N/8:R;TecVACf
8f?cbCZ4a<M7P_47KRF(R@O8L5PeU95cdARO3F5+BW+gHY]^D4):+K\5V6(cC;5E
(-0L,-3I@F#H2V#(>&Q#+>?V-HT(HECPgQ.T[J3F]XT^H+[1OT)EEba;cTZ>7d0B
KQ9c80gfLIN-ggXO\bP<A2DFY-<FYAH1K.YUI0NI/IQPB9feDOL:)BF#WFJ9^B=3
5E&X4[J8d^>THWdNSW2)KWYf.DCNH3+RHLEaX9-MJHX3_4#e)?4FOYV99KLD_,^L
\V1a_c?:EfA\f/Dg1EW?\P+#>:?Y;8T1@OKI^:e?@c=1^W11\g-8;UM<\&V2MOID
J=XNIS-/cAV_V8:geP#2=QX(43UC;a8bM]A/V[a[OF_J0-F)gNL_2+b0,F/=0O>F
EKFU,7<^\.Q_bP4;0F)-[02_R#S;IYZWggM/Fb]cIXJ1CZd6=H\Bb4e<)/?e_2OX
)dRX(aKYfP)DMBDfUf-HeX;Z[O:VGQSbU_UWV2EWR#N>fQR9a6gX(VV-E;=67Xbc
(3Z,+H/:-&-,M(\HNXa?>F]H&;6ee<G;cOgS:P999E6e_T_NW@?@3:J0>gGdGSIH
J)Q]VK?TY9#7PU+<=/b2LP,,_P)-K,&<][&PIEbI[E^e0:M;[Kb>@N(6Ff._\NL5
VUAP\WfAL7dOQ536bHQ-=@8-/126cGN52RFbWbNDIC4+S3a[S[X8A7ZHHMXYAdSE
B+@[J>@8RNQ7E]G)T6(6<M\(1&^OgPCZ?Ne55eIQ&@0AfXM?Fg#TW_N=AA]TDLS4
:gCNgJSEDPa\),ZVg_O(I6d<fdK.LWGNS;X8^7_-a624SZ.A0\-R8UFYfD>6cYI.
.8E4;MTb6EC?Aa7Qe:ReC2;PIF<;VgN8XO:62b573H_AfF<8G5T1-BcP@+Q&R:0T
>72aDJJ:7N(I?]<44--RS6M>e_dIUP[D-]0>C;CZ:&)A9SM];H]+)=^/M0K6C?1-
3(7Z[76M2dTK9aQ;[6T9]6=fW/F3U6-<..3J5>eOU::E9FJK691/c)a0F]=g4<KO
4DX_/;fCN\8M9-3?A7bK.JNU(=UBMd_g5^H^G)NQ-08P55UP.IK;\0-]+g#<X(XC
<GUXHRAM=?I-?O7RE#[VV,CB7QM\e0YDBN/70BD#]#_P^F+BA>ZW7RW?DK,_aC8<
G5\+#+UBEHU&92M;AZe<1KNdKL4-7Z)UacfK]V+F7KXLW]7c/-K]KGSf=Z6;FfO^
E;F_+dD;J]-7e-HH;0#(NaQ@DGA)]@-\aVTA:JN_>O9c@BCbM(>QIM.52DD3:Ye0
0/^<1>EZ9ca<&3^.cEV\g[Q49We#YLD^#;TC+XbcG_Fcf;:TA8.)+VfDH7^QO4M+
/D(&Y[Id4+^BbW6I&(ORd53[Y=:M?ZE?afD__+g;W]#]]?WY209.DBYQPD^B\ZDZ
II6^e]T@^:Q)2,D[LP>5DfNGLGQ^G&VfNV3Q&b;(58>])gIYW0Y3B=ATIJSD(V#F
:N];:3?d.9eTIPY0:X82XSf8;SD@S1R+M>IbBG=2Y94PGDB[d_.+/ZTN#T,SWPA]
WD\A6b^^/W]eOHRKTcQJ,I>_IZ_5JbXe-9V[?ET#YdB8N5],WZWAa[/><Hg[5X?=
#G+(E@>1f?c.dc@dC2E\ec<;NP,62^G,G+[bEgd0U[EdZXEIg2S6.MFdTC:J[>Bd
^&QZTU&>d6FV860\]?TM?d+]7(S@D[\L5e38D66/G;GE:2+bLc:EZD]Gg\.>,J@,
MecP:b)MF0VGGZH7ed132_,)a4-:FKLULM/c(5-DC^<WY^?bJ0Z&V\^Aa-_?S5ec
f;ZRb08VR@0(WcJVeY\Y9:88/7&Q-_gL:9Qe+?g8F<\Z,9cJ8_[X^(GCaN1##M.)
1EWgDEN\U,8fP;P+.Rd?Sa>R1R=0aTS./GG&3U^R:9_RI&=HONJd@>),5A<f.6AS
^E,7^_DeGPc<Dbg3BFUTW-b:P4\PII8]<65#<@J[ffM21E1?[N#@/IF&P>SIB^@7
1<9NdFFVdG5[Y:;>U1ZI/cFVc\A6T07IS#FUX>1f[TE^L)=[,0fM?W?FZ)#4NC;<
-f.5R#T-H[eITAF_CaQ>8LQH].Xg3eF[QBfed<ZTL20L_@7<cD&C1EEHY62Sb6OR
E1dfY9J^Wgg?FVCcN+]gYbD3#EXS5(?eUJ?-M,L2ZK_c&\fNN)OGGY(efa&-T-/#
Cg)VU,60\P_JY8A=-J44FXZP]+G1;TC6#\ce?g)MU/(->>I?MB5^ZJ7W#S\W;&E^
gW/K-0)K+L0N;S5P^Z<cNCLATU+[S>\OBJ0>LKWf6;4(d^_C^c=E=D\KP^20b8_-
E3>a\ZQSJMI0^b<\)=f2e)b0,JRERWOS)>CN)1Ng?(DSV3X7XeE4G)R=^TT--A&(
;aC^6+_eK_,R+ZN][IaSGT-M&98&MQOZYR\>++0d8CeMAA<fcLL(cA@RXI9a,e0F
FUBPW)6\^+5aPg;G9NO#-P[K-6>)d6.7@ESe6Yf??Bd@7:D]5(\#0BV]F0AK)aNE
<Q&FK9fA](GQTW#2/ZU6A[(R@\,e4,)5]]0/_9==EEG:U@C<&3QR;9OP.V&e?S=B
_QbF.54B?9H#KfabLXR)R2b,(=U@=NFBD=T\&\M_JbF6ge+B.3S4=,<FgDWT-CH#
D77<YNecO2A9I5X(843<,d(fFKVbC./0L#26Q.Q.8F:E(<^=(DCA&M51CY?E#H2b
.9XW3T?gI\\QVB#CJUGS73IV<_L4CO7aJ\5M?2R\VD&=R]9+H5U:N4IHdKgNf\EL
I]VRJM@@eMH79eDA+Q8PXHQG.ZA)U)T6.+VE[(OKRO\A9.P.S9F9-2^T&LVJ8?dX
STg?Q]M8)J6LK&MK<944PN(.[45O>[RBM+)>1]VBdHE8S;gN@R[JPf/IQ+_(\50<
=OJ?<V@TGWR@^9a:9^K^Z3B&fSM+=R0I/N;RDKTUZ[JcLGg#/<)BGBPLNbT3XHPF
8U#@38@/I+fGf\=.13G[@>TQ3f-K>Zc2@WQ6;QNP>a&@2F[@PHGOFP4g>3M-A;b3
=Za)P0UI(-T=@CGGQ8e;B8B(A<7ATAcN:<<4&YJ:g6Y2#a#;9S+,8[BJ?&gD51AG
\+EA1OC_6#V(&B=W(8CEWeLHSc=6,P?#<7B(T7CABG\4,PaR9_a3ZM+VO>?Vf]:Z
@O@W2Z@F9NW-3#\A?#E7HXYY50&;-BbDV.XT#/<WLgK]>TL(^g]VX;=(#9)],M,,
Yag<B-HW(\D?&5O<KT-+R\K@cI).1eY;.3Z=>[eI0)YXNWZ+EfK&D7;Db1VV=QK6
#^@QD7Z[#\6X^VNgL:8^1P>_T&3b3&TZW+3Qf[bf66?fQ1LAP\Q<b1/<.O#BfZBN
(J=VLE<Tc.8,>\3fG^O#QH4eYWG&+)eH5S,9&E0DEHe(YD?T^?\SZ=-=GdHN/T;?
S4DO8-<=7;[.OfU]VO35b53QR3>14D0DR;;OX6W5F,;28e3T/eb^1d43+7+.PJ#D
2H:_WFSeZTZ+>M_LK2,g=GA.N5ddIcU[(Ma]3Z/(A,YXG^bKbV;F?3;GFaE\La-8
U^W]U/EU+VT2CHeE?JT<.&SJV-H/#UaJA,+).8bg+)>^bKVe&a>)DCbRc.CTC?Ec
IZT.S,/H.1<,+f@N:<FC:R<]#eFX6E+GVJG7K\TH3b=Ig#?4O)9#WFO@KPU:/5[X
:6cGU0EP[P&/H\acET_4P_L=7)=<USd41DG3/A6)U/34B6F5#HH,8fVX3@I]QU32
6O4,3KGNGT3\PIJ7e9D\6[CW/Y#YbBU[dAY\?.fMb#3V_ER5N[7J7T]QbBdT?1/^
#JARO(<R=7H-0]43O<Ya/-YUfBP4_F:&E4X&gfM1f)<^YRZYNfd0;BUab65AF7.^
9(7LQec:+RX/KZZ1^F)41ePO7T[fN<,FQc^VeMPR,08C-OK:OFFDBQC>FcH<NdC?
F02)W+EU)0-4S]SS>IXWb\V9/UVD:#6_aJW<MN#2<IHWA79<8J8Xa9\aA<G0U,^P
;:)9#,g[a&eM6S+dR+77/EgHN:[T&JYLaIRB<YNLF8Y,3.;D8F2YCTS23YR4S)A<
1_[/-Q611Xd:B>7?ZZedKE=YU8GLcA^8.L\1]Ec1;.0+@>4T#-\HUOd5H[=DGJTS
#YJJ_Gd4gRMa>(g)Y&7&(;FaY1)L1WO3=1a7?WZHB-dN8RDEg49(7g8[;G8UHdM<
[HU-W;IKaIFZYE92^1RX0[TBcfFDM84eR92E4\&Z,SV)K^cc)O+WX[0S:)TB(Qc.
;/fZ]30V()1T4:.MZRVB&KN]BZ^<TCb:XR0O_-:IA6.&V]A].a?K166PD\J3N-0X
a8I+FQ;ZF#@O.@G_#e-c+M18d]8I8<@]bIgS.K\O+XDLX/3dT@R=AFg98V)NagV+
8.(d+_YWSEB5(+B?<FH4)@.K.)7K10a\AV2+XFFB)K3M-4DEQJQP+ScbScB_gea:
7,V9c&]b[fYNJRCBBdA1LSGTTIW^CUYAL;HcR0RGT3L;g4gM)a;1U#]=B8LCSG@I
IWGXKIV.0cHCW[NRX#E);ScB<5ZYH6GC/C]@8:a-g#6+XT?gf]QPCdK2PV@a^B5J
14EdF@fU/cG2)_7e(NM/_R>;D.;g<9Q?3DN63dee8D8JBT:.D-=A];:(ASeHG@BX
5IcdT.:g1Z5dPCLdQdaG-24WfbAgdaB/H,+8RN]W-0L^TWB@V];MF0HGfTaW2N2K
IKeLBLM>K(;:VX^EWfUf+5S&E-Z,2f;2&4:e/1V^^RU^/#KBaEg@@eG)eQ&R:L=Q
7^Ka<]=__PD?cPe.S9:2D>,g^FC^36aaC0C.PT)A#]Rg](Jc.D/1MgXde=V-8M68
<+ER@U1=;T^QDB0-+Q8[WMIa>&E,:89cNB-R-CK>23J>Cgc)W_\2GYQPMLWD6I1C
A;;5bc^CTC)LGMK\0cO3IBR5RV8D@X4[0gTOaT2-G]YV:#9.#1C<2K_+4;dD=G[V
PIG#agCG&SgA[A)Of:(H:/J(A8DPaU4>LB)KLFRb4&KB=XS>OH\X51B(]TYVfeCb
9#4GGdF>]e//?gOT7A-+8J8OLG&N2DP]\VM5[?7P,)e@NDJ?4ITB9U4OO<;=B7+?
V[O3?VN33WZUD7P8O;ST7D3&.f#;,0[(/g1fF>]8.aUS7e5MLCKgKd7f6-DTO/1g
e-BO8cY4)NgKSFcR6_ER3C_F][MO=D0+Q;B?R-I8\g^6P2Db2]RV,=9[)V@PdPb6
\Z98EZ+HfJg>NB2,\BBXEWGT(SJN5UQSHe_@HVcTY@N-FY((BD]8I^M]+XF0Ee.L
/;bUWF:.0NOH5-5L-V[C-Y(092dPW8RA#UQD(F(8<_J1(aJRVd_I9>e?#PMgLJd[
=I#_<RM)+Zg?Y6gWY?H9TOZ4EY+aKEZ8.9g^\8;Q3,?QM\JCBYDD:J0f>_]gcV9>
(dLE-8HcL)D,Q(/97Pd^bH>;S#f<Y5YS>ZDUgQTO5CX8eG(&@fOZEPQB3gU8cTO<
^/-1PMU7H:+0OQLX&.)#cY,3PbR0=?I^J=WYWb?2P0DB?&Y,NO_.^TPaFKKDK2#R
ca,BA^c\O+WNX05]9QI5B=^PCY8_O_0,dO(a[bA9@^F@-T-/BDf4S1T^&>e?]9B<
bceIga>POe7@a745g(UF(A]78DVD76+/KbT@QTA>ZGd#<(/;@9J7aRR3S[R3,R:V
,,:L6]_BYE^70P.fLTXN&]FXe/^,b=AE/)I\K4N:K(b<U\HF(@Z;V<E5PPCS]WF#
#\H=[<8b&X4GF^ER4>:)S8fNUBCZ5(F87VM1KR<D43Hc2a9LRPAE=H4-YUZB?CDE
58QPQXH]b=\C+1J.KQ()^7dcSSTQ\^@),P]3#A@Q]?/#\XH[c2&1H+-cJ_8^I/=D
-)G,4P4O:EVC4,3C7M+JYd-T-WU1Le?0EK/Ga]b9dDM9VfDS#I&A^:Ab?GJ6S\7P
^T2G6Kd1P;F?71##\@57JD[,-W5O+GX?f3-\e<<_V1D7RWPX.]dJA#-Y#_:#KVYK
aO^9AHO5-Z1eOCG-X]AZG0..,CQ;bZKdQHJT/)aVCW?/H.[ZfQCf/1O[D21_IV-=
aSI9;RJ9cI?^.9D004b;H@06g?TgE:UN]-e\<7O_F^\FAOY1U7LN9Q)C<91>2?<a
F(PV8)]?TELGa,>#[VU.RQ5eQ04<6YGMU5bJJ89=Q0P\;L/N\VI]A(5V_ZB(C?aL
,C(^_\XUO]AHUH>K@V_F1AON_?/WIM?C-N^^FbJFWBbbPed/V<53I/;UK<(?/dDA
R]B.RO2MV]Q\RL_G197<@.Z.b_Sg-gg-[C6I2(<_5XJfUAA/.U8G;c^]X1LT6C;3
?bF(=gee&+T0P6>\&A[<I5C4W@JM9ZEaAK/6&\d8f4MIKHg3H=A2/2K_Q--(.0W8
X;6D>Q-T.E=9dB682V-OCTMG\VE,TBLX0QYJ6XPKQA\O=AHNYV;gI<W<e_7F>@ff
4J(1ac?Gb)DAX0&>@<Z:D[Q>HO(-bT[.YH&FI/+JF-b1[3^_7KTQ2W,92X0R9^J.
?N]8HfNRU0WY1:\7&M&HPX?+,+:&Z;GJOMV_;A[_E=<eZC;N0Ig89.@d-?,5Zde?
I&eL],/&1GG/BX>:a?aS]2.1>6C0M&?MF,Q(;JfOVbSV#PZ8,Vc3&T&O+O62;SV#
f)EBcI)@,[E<daA2V#a/3RcM/-b@fVQ&WQd?32B:Ya\UDW>#Vd32WcE.,5?)QH2a
9:gA?A7Ca-f\.3==9g-BERde>a1a+R-Pe9S]5(N8A3W#fFF_V:^^Q=KFD#bI^-g#
-+J&MF-(gGPI/@:+])Gdd,-#1-1:&+VCV?82)[OUUUc6D8JE(?K/=5YT(bG/ODFK
X)TC<E=KRHW0OM/B?[T\2NU3,0-Lef3BWZO8<5\g=R_VG0bbKZT\EN-EV^=WX-aA
CW#5>VIS#ZZ&1:YY/F?]3d4-9/+A>MY2#VVP_C#LNZUU(Y\0=TA.?]31YN\5eA\V
?Y9+#cU=BP&B7L=Y=g;gTI,eB/g:E>.W[@/ZG/1AS>?S@KKYec?&<2D3T+R9c=bP
V=;geg1FD#9,B;LMQ./<[S=)=T[QP&:4+Y1@DQ^HEFJ1XUL,T3gc<fL0LCAD\9B]
GILMI?^GS:;AeN--.:P6WcR3<;Fb,_@ReX9ZD\8)2ERP?&=b4A[Jc.5P0Hg^4<_G
-&0/MV3,X4L4?aMAJDfa:]9/0^[Og4GK,g7VAHIDU<JfO&NV-5ZC^8X^YOYg=5>(
F)<7F<N;KX97Mb+eM]:D&1;PMWUHI&.UXPTaA_6(-_^;5I<@cQXX<fY+X&[^+_#A
=Kf)()3QL&^Hg-K(SJ#&3Z)dgSFXW/4F(GKbeFTQ?0OO.8d2b?4cBLUEH;dM3P8Q
\@,Q31=6@F[T?7KQQGPT^>_-MEeP^BO?6C:=K._4e^HMI@MQR4XK5d/<f(-\DdGF
S-,5UGf@G5RPTRNG+Rec).P2(V2/7+LV[2GI-\T_;M]VMI(NJA:FB>QbZ#IR9784
)WSP]2W@EQG(0CbM3&9JNcN:(CcFYKWf>(#-T5_M>SAZXbQZB.2<KJDd3Ege23Y\
A@_b2ccAfHVPM7?5M_D7b;aeb=@RY&)#QE3Ud(5\X)N6aEFZfDgCYRWT_K:af+@4
?7R,+7466B1D4-=W^J5<W8Z9gg^<SI8XYBZ=b;.2?QaEbI#=FVPLXV,De_:gTX=1
g5f<5a=L?&/d6f77?H0UA)Ze+>YB[AYZB\Z>K2(+?GWF>^327L)+Q?W>LM=D+_1E
V\:7G^HgO&ZG,TeEfSTA0=V6_8LE_EDQ-F_(J-[TBP.Yb#Z(_L\^f,,ODTZ2==f;
KWQKA+N&W-05(,G2aH-ZO40+;AW55c4c:U^X)B2,.V<+G,YK>-K/7)#a5?D/K9]L
?,HcBN66B>4\_N;#.aIec9(_T/O7S#I81P+GNE^I1:R-)=-eA#^]C^MR:YB<+332
,HQ68+GMa/GI.[3@1GQVJOJBQR5.P^>L3LKV(TW.>aP^9VVS[N:E&^g[,?50.[E)
,:-C;J]R,#3@XSTaP6O)-RUYTMcH=).FPM\e<S7M4<H/>5N;<4.=@fcAURR]1XB;
XPNS@CRK(_<Y(>U\/NX-984O;ZY0GO/e/QL>:CQJS/1g5M=&J&;YS(c/KL+01JfI
7_6NJ>7X4-50P.<UQDR&[1^XQ7f3Wa@-XKGN0=a5\Hc0(DfXcc8f3aJ+0U:?;&&Z
d]6LH6DK<)JWPRUc9XWG9<NX4a7\@?1]eU#UD?(a.[P?+7K6QW.:IG8XZJ]78cfe
(3YC>1,WWSg;S\DX^(3QgV#W2K@L]g\TbB5104NVaPcA0Z[)+E+52Jb\&>Hb37/E
2PEX?SQC9S^\0A<<.>\cNf.92=>d?3]MGHfT5&@8IR(Kd(NdBEf:c::/MKR#1WH:
71Kg0+@1eQ,#/H(709OLdLX=O.L+6\d_Q[FTG+ZWYX=6;SaMc>][R1^SfZ0E:EUJ
MHPDDK7OK_4>.D3?(/1Q.W:.\)9N)_X##O0[2e6WS1@XBH+GR9E9S6<]UZd8FaU2
(b:8Wc-6ZO>eXQ=:X:GX.)30\O.Bd-<7W+K8[HJ)0++EaUHOOXP/@)UG]c3(CcS)
@#d1-aHbd9K1Vb+F\(P<A8/>BWOK^M6f2g.SN&;a_+_24bHOTRH(-+eU0@GMDNUR
9CTS0N^NfAWJAKTA]8_OUDNb+,5YXMAJd\DF3._g3OX1+>LRY^Y[IYA?G0\2Va#/
\(g2/WE0FJ+-T<e8,4TVaKGBCXFL6BLKZ0_/(88KOOTfOL9[44>#6J[+\11.@fW\
J17]K66)1.3S[XY\YB/=S5+?Jg1TFN_JR.TX<OJOG=f3gQNETR#5c8MV)gOW[Z0=
OXbE5KSLGNZYTI[\WW1B6>,.^8<_P.6Y@U)Fab-G=b,KcQ+PKH3Z4,1(VZ5N?@?0
.G@/.C9XEOA0fCc7&2+1F:MW-9_-9G=/RGg2,/ZPI<KWX&f3[<1VC_W9XM(_7b@e
R)1ZM,/W_-GLU#SIaG^71@#HH93e.GAOSOW]9@<(5fF-?9JRd<_(1M>==5&LU7.C
dI8+XLPeC9JAH#ggZM183d;PP\Q_TPS=H/T#-AGA7EN5]9Kf/;\8/XRSYA?-TaMH
B\E3/97TG99I3LCbe6EXK\;3f3dMWSX](=cT_M(f?cLN(4/I>W=&O=R4.GSURP15
Q<UCLbZ-PCXU80EH_I\9Q/?e_Fe-&KGK/Z+)2K2ZCMW?&7J0CKf9]H^--VXc@(_<
[T\7V5Ga_/4PX_-[W@P?V[W6T9/[IO5P@>e9F8IT5eQ;ZdK\66/e>?19<14QFTfa
fX:G.ZU/LYZAgd)VZ_?:W]>-OGJC+,-;a8S.WaB_&7H4?M&3TD]9;ZUY593M>>N_
.gedQ;CR)&db,@(7+RBfeB88)5.(ZWgR8YfA_M99EF,cCgM&UH6[,Zf520VTX;1L
=@B-,8WWO?C=L/6;Ebb;:D<Af]\HBJ4S2fg=XS9O(\RP.f[FS0fBI\/4LI:BA]0,
V?d@X96bW9?WDf3a^UK<,F[9@<d/O5D/JW\&KQ^#/-,)@.R@^;gPg892Xad5JD<<
=LKB^02]Ce8G??F?dV+LbL(6M(PL@VG6\Y)TD;3gS7\MI>D5@cC3KV8\4)abCPV(
(#XaMc&,LNAPf-C>)0]eI_ZBQ]UJIF2M@Sg4Ldb\aFgfK/FLE,A8K;877cZ2A>MX
A;^=IAJJ1AU\EF<aKIL<E^-=<CLL=7eH@:++UKZP&GJ\5d=dM=_J+UAfSK&)=K#Z
MVe-#,+D/34T:S:M3)9O-UU@+=75#CCRaQ\BF-;+=18bgGOVVfaM,^H\&KL_-Zg5
d1)d3<V4,.WOeP_CL@:3\0;SDD;FS+d0^>GY+5HTV4=dQP20HMN5]K+9+\<9aXMX
8+2DHA&W+QV.#62B4BfY@0;33f5aO9a>XH5_(\g<KB7-U2,MPN:7aUJ&FXa]NG-5
NQ0.ZOcUf52H:cD\NGA)E?dK]X(Y/NBYADffVJ/T0DG(MYT(^PJB8H2S1CAKKTJH
W&?</H,eI:D:a=)8NN[Ha/Zd.)0KW=M;IBMD?Hf@RV+[F<[2IM9)LB<=Ba8OcV[Y
3[=?2WX8XS+HXH>Y>Uef\[7S>0:S1c,<-0b.3M3^/^+P+>Ad8T5(--U[>JW[>JF3
fD1U27cBIb?1;<]=dCSY8Sd[:b4FT7EB8\ZS.8bF1A(02G.SaBYI:O&Md^\\SAeC
&F08TOD_WKI1dQ8([].C[=(cB1Y7TH:RAfS>E)P^\):=]^^ENJ+ADNK/=K@_3T37
]Y>.a7[X>)TC.;bJ7]4=P:NG<];A6V:[ICE,-R>YN3@U-\V#?8dad[:>]:0D3WK;
U?d/QR57C92,Q>Y7WYYL\2e[(?:aY^?7Y./Ld0^@@I98H]=\WMW/d#g:\VA6TUeM
?E=4B\Pc?T-dAV6SMRZ<^,4IaK14a5/b@Q[bCTd.)a?(V)YW/5UH@V=dAGQ7C3W1
/>LWQg25bPd@=DY.>Uc\_a0ISL:P((UZM83Qf1]R^K&Ea(X]_/DU0S=bAX68SeC9
S^Ra.(f)#J8+IWc_[V[=MC7@(H^.71&/E0=NMW:4Y\cQTLWgS9H[Q,[2U,=7>eE/
098=8@6BZ(aT[V9/Y(B?MBd9Q9JdFNb-Y.JW]fI#J>A\G6E(YPbYce[F_>F2VTP8
Wb?<9gbgT7+(/333W5FTbBE9(76.]DF]eM:&)^.d#QagYQTY+TSPM)03.^,VQYSX
DG]<7Z>>Ld\Q=ZMX,+A[W1UcQ3eX=7U3?/KJa]M1egFK.H]BR+<RBSXQ6@/4O73A
eGT#\WJ?)X9gL,78Y;28OP.AZ+EW#FX=Pd_><YHcc@3f/HK@<T7ZcWf[X<,11G7/
JGL8[YfGK5I-HbWR.gcW1f[eEPdD-[V[K4DfM46]KcddY_+66Ie)2IG^f^]56@(\
QOU:WJ=\Za:+a6fEO4TX;&5bfLU-^J&cdMQOAE)Eb)]d<HPYV7XJTAWCBe6IJGgN
XCHISWBRHZ]LY#_10@ea/)9bbWT9(J92QgUD;5IR7#JK1:UY@)9NQ[WPF[J=Xg9g
13^9OIQ+C4JfPY+]bXf6+bMUf]C#P,+I5Y,]QJD]:7[NO6:VEf<5?.WO7)H&T>0U
R-]/=X5#<ZLD=.f.\OV.@cI<>FN+&=VcPQ7)8<(b(H6UDM;M<fQJRPU@7@G_#VVe
\P<L7B1dVgY=)3#_#@f(SY=cD8HLXMcX/638&0#Q?ZeGc=dP)YG4a)ScQ@>S>44\
2<##Oc=L4+^^[T384d;E.E@GQ<>SDO&@@0@=^E)XYM37a9C/JN4E)41[a@2Z<Z+T
7PUFaW9MV948g)HcPH+U8]7ONK-U]1OPJ6\6[e0;)@cL2>4MZ4-A&\^43.(X[@;\
E/]SCM1[gD4,fMNULRT^SW@a+aLFXAL_g-I1+gBG]RCW4_]2Vc:;/LO8]?[4;XS9
_9fU1SB0&M@4?N6S6;&CZA@:_U/Bb]8aZV=YgffXC7P=.K(ZfTUA7B#@)cUG#5(b
>)bg<HX&S#=N7>Q35PZTbRNE7K8@<EcS0)b<?.>DL]).>/ZgcDeN29ZNAB)10#dU
GN,\RHUX8\YMd8LX:O8;+=;7F\T/9gHD\Q#/<Ef:PJSWa0]+HG5/gJ[&^8TL63R[
=Z93^@15W)F3B2#3;V7Ga@=WWDWA6QGHJf#W;bRa3DP)CJOR7@<,X?4RW11O;/CP
Mf4+HUece>CZ_4VX1UZO@]7G=b4Ne^TT1)][cdJLb>_/IDcN\K>bbA)1N->fD[eH
::&#V/Ya,ZPWFEW-\G8;[J.:Y\7O[[J[,09+?28X0Me&B4>8_^;WOAB&3HSPR(.[
;-<5.B?K7J>_S<>/1RRDV.Fg^MB2R5+(Kef>GOUd:YTHY7S.+3&>1[QgMd;g.Q,M
0g9[c(G71^>XB<18;7\;_63gWS5.67J7U:TUaRB);1#WMLb7#C>A[=?IF#PPWgCQ
gCDI1-?2eX?1OJXL0/JK_f/N7>AVJgg1[ONOR:d08P:P2@->DgVOK^E),MBN[@D.
E9DW[.8H\(?M/6W::ZND\Z,ST[S&;^7DG/.<?J.L.3]&+Y<@?/ST/7cICCE[3LHd
N.GcKT^P\-fD;bO)ZaCeMU5H+AgALFbT&O;LGa#(QA:;,;JL]#:LMT-.M<egG-]H
\UJ^ffD[D4SL4&g7MAD2H3e,)U[>ZS,X.8:<K-XaX3f^fMAH]C,Yb(M\M]E#Fa9@
Je=5+FcDJMY5G:acSOd:b\VdZOb8d\X\SdEf5#M.EPf98H&<XF6Fa\E#2MP4IdMB
PSZO+VEQ3_W;<P7b&R92+C71CI#,E+?=e7D?B75(Y-a>&Hf\<?R9Z>T3Z^I;3D70
IJXN#\B(g9(X<9g+)D>b973I^F1IQ13ZTB5D(f52F/H6+4CDd7ETf5.@P=@QDc#?
1.7e.I>Nc2OX[N[b?5)&D2&R.D+JBV<eGDaG#8c)H]a3UU-H12SBNTa^RfKBeO+S
A+-3(X.&?&KBTY>+3^@MIAIAYXE-L?NXONE-F@:MP2:-#5;4T.Pb]f,\@?K^1]GC
O0gAH)C[eE]S\0fGe:cf5_EE>^UL\1D6_d^H[R@^K)5XP8dPY>Be:C][F5[Z90KU
GZ7e_6a1;dHU5)(,=gWKQM&EHUa7Y^3G;^,-fT]0@F<T1]N9-_7)[V^SYRP.TD:g
0f.8PfZW-gOCF\dMZ3(TS0RYUEb95a5YEW]T]R^YagRNO2A9=^/HS1:D463GO(PV
,MB-+,?K5)Rc-MT8eGE[?GCf72FYefF0H=Ob7CEg0M)PZ.?JVS2dc0XS2U14CRb4
RUD+L[IN#<I^Bc:U#+EYB@T=45-@e:+US&^?906C<8T87+g2S);?,=R<L,D>\cKg
ZH0V<NJ]_L]acI><LY8d&f/VX[5ab92Kd5K1RCN@Xe-DSaf(BS\Rd65CG4FXPD-L
\]Jc^1JgYV^Z>,6_O;9W;<g]I\NRJBPQCHOSP3cD\A93P()HE79];BG@b03<Z&?I
f]65aYN+6UR0BW8.IfT6QS+-ABbCP&HTI46>G[?9;g;1b^<K<J/^?H.ZW)Y=C3JZ
45=5KF7G(XWL^F0T??8F2CORYa-[LUMQBb+fF-OP[AP]FWgAJ_feMZDR#4.+fHF&
^09HBM9UVC>PBGMY@Ad2Y^-.>?cHG4/_.>Q2F66&UEVZPFN9A5S9B>ZR0g+X<G.f
1@G&)H2MJPT3cC=KJ+VdZ01&,]0YC\;H;&1FSYIY:Z1fc/>HMVF/QBA&\-812I_,
8E_^]e8:aG&a?XAFP6-=9>Z<:=3YJ3J94XgT9&Z_YffTI)55CQ_?)<0E\Q[()[]8
V=Ja_ag&TD05MF.SJC#20IAHA(6[4/FY\5TOYQ-C7\ITVg:PFE8UAPK3DKEC5#d]
a139<U-WfIY>FC8EFWLObPga,Qe.[KF+CdcV6^dU(((Me^PUZ#NEH<eYdZMS]dIA
M;57-Ud>_;CcWBTgb<S+NgG7)V[DBaFED.=2a^@1YJFc-@4L>>\g:^9MZ.Eg@ce#
E#KQTURCJ+V[GWPZee?]BMgN/B@?e8^[#&_)B\eZ<CG.F<cec=Xe6)bReGA2FbL_
;5[EC)]:Vf=(3(K-Z<AT3VW9P&2>],)IAP;;L#^CV&bBQD7\H_HL]LaGM^8TUdM)
Q6M9MQ=FC99M6:E)D2.KHRL]KYcKEWgd_,-N^]D.K-\..>ZCCVFZ/J67M))DJ>:K
_RJR57aGE.86-275d&XEDKTMbScW[&VUdb1NQ[>X03;d\?=8U=X=TT#K/>\5E6G:
E>1J2?Gcg_9:aQ5YI&?cJMLA>)?c6GD((5f=7G/QM#2RAC/CUMB5+b&T&H7974]:
E,?+Z#JOQPKNfI30Wf6N=LaK64dY>JKYUgZc4PO#U)cI.[bH4-X[2eSI(F4>C&P3
&U\-ELM=NcVYP9,;U:9FS<-8aO?XP):C4JH1LW6;7KQ;2R38L3]GfEFZK<Hf<?JL
QE5105_0Q+/2=8-fGPYJ4T^cRXNV#&Eda7\&@..)\(MYX;YO6^We=;R<^]@]@5g)
S1U_8;+NI1_3EB0d#3N4Q8&f[;L@,=UJ4&S6IY^;=e\b4d72#Ad.f?1CE<FFA>dc
IA-gXK,F[1M1bGBc>FB=R3@?SA4Ve^PVC84gZ57Y/]TU>=16E@97>bW>#+@86CPH
ZOS:I:&-@_4A-2,1=ELB<;SfRg:TgN]8_CXC]I,.3J[AbTM^H2(-g>0XJKS]bKYb
;.d7W58OG(dMIO<AH,@J^^E30,]P_#8<8aXD0N0],L#OD_ZbM,<AUgX+&;2U)3&Z
CP.T9E^QQca\[Y&4g(TE<bQIWbOXNEF.\9YMO267,bP?]_=\cJ5fU6W_;I-TLWDM
a0PL0YKg<:A35^:QG-=_12_S#^9>cU6&G1C#^9\B+X)F.013W+d1_3[FB(HJ1?b\
NJd:J^eQgP<;K.2aH8CYf)(UZ2>R^gL^U)/5GRFRS:Q01ID?-YZ-(J_DSI(2->QL
S,f/M]&<XLW^gf7\O]cGGAd:UC14W<[@#T)PK(.fCZ,cb]<YbeM>YHL#5L9C_W[Y
/gVG2ETA_10UC^GG,S27X?#I,8O7IL@Fe1[0&7SKO3-1MHL-7ZW2Z[K>JU_-8,@S
_.#Xgc:cGY0J(_C^VM5+e<Q6#-X-7O4Z[CH7JF[&91@T3X.&+JI\Df46c;2)R-]6
WdK@B-cN]L@FG5/SOf0C9f2O8cY,8R8E8KCSXZT7Q=W86S/\H.8Q4N^=XME(IPLY
IPX9AcLB\_V3cWMBHQUEK>PTXKXKa/eLFe([CX5I@b&Bb6>1I/Y&6P[0<b##9-R]
@_dF8MU4Ua>Db9Q+(M@)1X7OZ>0^gNgGUgLgdBOZ)Uc7CZ5g<1/[937Ff_#H0V_(
-UJFE]e_?4@XfRH>[c_:d]9Y3+f0\+,J)Dfd:&NYFgM-83Vb[_]L&96C>4fWK;V+
>\;d2U:&K[Y3]:W5[K(24a&Y^K0C1N:6WZ3IZ34Y^?aMD8+?\IAPX+L500;d5:F0
UMS_bN5faIT>&FP>Q#N?+^3/.,3<X7g4L@Qf)0SLYL-TAU0<Ne.I5VA8E2N=;PKI
eQC<H3c00a@=;:]_?[7@Zd_9.=LHPE4N#Ug5^W=IIR8>CU@[#S6GF0^2M(#ZGNT)
f<WYRL52I[[X,UH_\V;R2;c#e&#.VP+YZ3X+)HGc;NL9d^/DK\P)[<LZ_LR^X:1,
fR\fTBWQAV-?L]CJ=c:N]TOZPC=ABE4@+WP]M+I5&+?W36H:Q]3J7P>e7=4&faMT
=g2;]M8gC6BC;1CGf)Fcf_WI^4EPGY,g4-DcFC+X4e_8JR]KG3W?GK^FK0@CeK/7
A>=>1+I8;2DQMcF_OCg?VYQ668,/Ra0eagEb\;\Sgb;((SC\I^(@?IH&3a&KLgg7
L<e6g]c#H>4-QV7<XO/C[3-[6:_)_4\;P.eg@C:4[^QM3VaO(@a\27QX;4OO?V<4
L][-bT)#F>M1^)JAg/f:CQ7O^--:JA056&2A<E[B71Va&5Q4K\^_D#OZ^H[adXAM
A5E=I(=&V\L@D+5;RLYD<Wd8/,dP./A\2Od71D7_1>L;eA^c7.B]XI1+P;YLBF=F
>B.a>\;Y\3<2\0:B8Zdg?K>\0UfK2(&M73X2f/(T&O(7:C,BH;@\Bf_H7C5?PG@E
/QLMTA+)?;a(-YRT58/Dg+?3QB#;8HF-8A-,P_R7_]a7B?P,;9f93K3Y1dEDL;^E
?Je3IaeT/3Z:E/P68-^(dSO#6U@B0>gYc=e=DTfE<38+eI84N2N-X>+R7]B)?Q-?
=e-?_-#:)4+Xe;:6F=A)bF</.AD\[:g-L4M409e&194\8gGF?#E]a[1T]0WOYc]d
#?H:#9=@,?DQB.9G4RA<CLH^b6-O/:]VK18HKd2OTWXd3I>&eL)aVHZVN[HY7<G0
f@5W,@U4]K.3]1D>.ZA[K],3AK2c+75^:X_9C227_Q1OCb6aYe@#-^T-<>Cc<L^2
?UTB29D:E;\KK@19e;09;fE<,^WI\?egb3P0OgAPd[#(AH(V@PK?Q?L3&d&_(ZJX
AQOJW-K+<J#-]\AJ[ZSN?(dDR^NDM#J9-EJSc;PSe8[BY;S?_Z44e9_Yb-f&Z4c_
X>HaeXRYA+K;OB:fWXaL6DQP0D:?_&AOB3KV\K<R?LEN[HZ1]OD^2@9CTR.D6<+(
GUVF),I^Y::RZ1-E.cG097\1&R4@Q^&#F/#^V\,<YLM1.Cda;gBZCWb4]2fWQ&NZ
1,[O?f_TCE1c@[BI&=(A^N-a/a0G1E_C>OO^93,()P-P^+L8G6I>,/Q@,5LA<>Wa
K#EcBbO,a3]]@[6^89#PA-8#,PX(.+3JDO3MG>3I0=1?G7#Ag36Mb7B?H#@7]<0E
/c\W\7<5Y)71PMI7Q1V[V],H&A1;IdbZ+5f?]c1XNF?S?QVWERbYO<1OdBdU=5-b
fgG)@GTV1C&eM\U]2,3UELJK0BJN>a?7(RN/cUcA1?cf^&C(=@E.:QP))d2=QO=>
dOF.Q<;2/<&9SKN0OHU&Q691>5LC<^Q\QQF).CGKY8SQf=gdg8]/:[gf/8V&=V6J
_eB4H/e;N\?KMG0MbZ@3EJ<:O0@\\3@?KGSYA_481b\QB$
`endprotected
endmodule


