`ifdef RTL
    `define CYCLE_TIME 40.0
`endif
`ifdef GATE
    `define CYCLE_TIME 40.0
`endif

`include "../00_TESTBED/pseudo_DRAM.v"
`include "../00_TESTBED/pseudo_SD.v"

module PATTERN
`protected
81+MWC80.TFDc-H^DWBe6G641_P1DS?H4TG<_dBC-HJWPA]Zg&gT1)WK@#Ee2]d2
R4=e:O2DU2a/HW+FQ53&KJQfG.<U>&LdH_GSb:JX7DcE++;L.a6+4A9MfZR=MQdV
+606[HZ80:Z>6(]VbZSI_)5^e(UUDg-Y:Kc3g(S3.^2fP,\-;(P?ff/<N87[W3+W
86Fdc^:^2,-S2:YEVKL[?@,^BHM_<\gE3>Yf_@8^HWB6MdWRXfN9LJD\8V8a>b-:
^(.5RQE2d,VS,_OR<@WI78OY.3DeA2&S1#[[;X-3T]LKQ7e01g\I[PNdIf+OP/O.
)gY=9We4gXaE@[\J5W6,FRXc_<5LT]bEB^J,@OAAD?:J2V-1g@7g_GDKEe3/NH8U
?4=]DRd2g#124G?(e::AA2>>fT1IAC7C]S,_9AE1VNB^aMX^_DcVOSd_E]6AH6VT
?bd,_Q3E,).QR(6FMQ^)A<>UL?L(fLR37R)0HH=G&7eMVX25/01]K+)E0_,9_4Z3
R^#GWS54Sb031RTSX5Y@P09=JM7&[16&6^>bGcJPEUP+3R&7Z.U]0)cZLde>).Yb
7ZY,;f.HHZ/4.IgR26GA3#N2B[,,>,C3KRMM,adXf.]0-5QPg=B-@>AI0?F>WPU6
P#/)0D0^T[=>)+0D@FR=)@^<LOc7)7N0K^DK)?FP:@4NWVFG?1A&B8a^a--97<>S
AB,4gNG0W7d\G(e-4+b^UAeE9NEKd\MSc-Z0YH10?<6[FX9bF;a2,Y=3MU=\eSQO
VV<2E[Md/.X]C[gDK?]YIFdb+5C9LD_MEGVN@EgLU@C;W)(V437db6W=-b+J+Rf\
+L[V2EaB3;GWd\3:8IW^=>]V?=/,?)U\&_(JfKF1?B@&LUZ)AUDRV>b9c0&B.V:/
fd<?6QR00Pa_f0222YO;#SfD[d.F_PZ4;aY#\</_ZHg.2bBXZ89/YGf#Z8=gB.EO
+FbT3AAQ82\N/d\[^]SO.ML]K@#97VVZPb;)2D07EK[.c46HHe2V1L#QFT#;1H<5
O^^^^M^1U_YC++^J+<#/P]bZEA)SDEX.NW^bRUS&K6?d8/a0:CNf_agXZXUg/BL?
Bf2Cf;^=S(FMb3F.>d+LJ;[HWPBCZ+OV1IUT4(SB+4ec<-?)aI=S8^@W:\T+68FY
e<GJe30Q][(CJL3JN2=fJM>)L;M-+YFISIE\Z;Y7)UJ>3.(.=)_Le9J/+-Nca?F+
/H+@g^&8;X_)J^b9FUWR?/_]>^,^Nf<d7_JDBWEI8TOeP+624FEF(WL^WX5>0&d(
U2GJ/OcI=1_ILUPHW0P]e\<VQ]/3M8\(,)W=^B,-GEV#^;1\=2LH-aNe+Z=3?34;
QeVd#e;](4T/He3QLbZcDR[\KS_(@V-Y2FT7W[3F\Y+#()F.0Wb-HJKFMg+S[8UH
O#@V4ZLV@D8(K[K?L#=D0e[?9^?>FegSQ]<F6dD3A?Y?,c?L8L(8(ZGH<RZ69>?K
LdY(RVHGJABb.c[JaE\U6Qe/CBD9CGeOGY;:MWPbRP^aS+F\>dWGB?AbS;JS5E]U
#PJB,+3C_8Ya^f#g_[RU/R5T+X:K_N0Y05A>=N,R]0:=BOUW3F(Cg@a)SC,P3CBN
A[;8QZ)e51TA5_=e;0O73NR_NdE^GY\_^P;/fPD<?dZ8D-=2DaO5aW:97RF3#J1Q
KcABK\+GMI^Bc0@^@5edd)A>QE9;QLZ,AF3@R@1JS1FP=K6ca2e4XA>HdC&\X9a?
\P8g+Q<BNX?HVHM4?6H#ORIDdceAUR-]SO(1)/M&.@.NZP(/[XF>BYcF>1E)0_RB
8R8:+V26SE&PB3b5GJPOJ&PZZR9:.+-<AANCgdG:b3:fDZ1#)&cMGCHV+d<<UgM;
7R7V#e_bYM&KOReG&7-f1&V7#[]Y<=P)&c^J@A,O4d^CT-2P&+U(\/C=bNaUV3K[
U1F/Q=gJE>+&U2TAfWGL>M)Y\,N7@.0BI(_gDQS\:O>@^[eEO6:[]BbF.d8,M3aI
dQOS?\dP_M:/a^b:R_aedM5[DD4C]RQ_f:]__3X2Q86:16?8YC[Q)fdMg\G7/7aa
3(A:Z3;+Y[V=^=(eBD2/YI9?\\<1S6W3gI@ZP=3+&C(;b-X4FANg7<eLLd[\]GeW
d+M]HG^KAT\fHIQ(,NHHY7];,Ed3KV1VQ?22WQ4OQB8dUSH/VXJ/2>HA;gK.GAP,
eQSF/-_PcWDe?0DA_/IA@bIIeAe?cB)K51HKS<V>CV)Y2LXKe\5//A=GQ=^(1Y?K
H(6g-+R)ZLD;ONPN_e,Be2[>P&9VRc]S9_01U/fJD=>B3-B5++[,-4@8(>0/+\D<
URQc5,TU3ZU^.\W\CC\.^2A@:3ML92RgT68U]4AJ]#:^e=GfFWHVH3dIO2,Zd07L
+bJWL-D7OQ]U9/dHQ\)WEL1C7JB^^S<>+SJC(_gg?Y.XJDRSO<P]4g<D/<;^>9#H
ON[d69QXS-F0)d&5H?@YX;39.NXTN)831I2^L;_eMc<(]5MSAQD+)T&2+_[g&DeK
K;QWWN5e3K\MbR25K;0(M5N>AJf#?MU<HC:[@SQ,X7AL.AcV]<,?,5)2N:2d1EfK
NDZ=0-R2,dN_EV[/?DF\NNZ]#JX\2?b7WRf-,0T/=S<Adc9bXf;LWFSCA:O:Y)4&
+cb9W?C\0,#PCR9,_Z0=Ta95)XCDK;gZ<6Q\[Q\R>XHa60=(Z?RC&:IbQ:MX]<@=
c[S^>>d#bF1&MB6Q&8e;B+CY&.ZfbT=Q8SFK1>+LYP@HB#AUEg-caT@5SJ(7?[fT
J+_-I+#LX&HU[7O[OHHLKJ4a\R+QL>UXaY736WK?a>b9-gaS7VSL-KD+EBY&0WOI
WLWfDc1fFEdBSeg4#)LY4LP9<g4#e#E4?UgE@6E@1eT;UN/>Xc<(K18(efLZ]62D
F^EV0Uf]F=BV\1U.A#-\<I:RF5>UB4P?1d8VV-I/4\7R2d<M0/8+NO<Z2H)610>_
2C?4LZ^.<f=^)N/](,\]7:3HJD(d8QL6_/KT#bMW-<#M<BRD=<EBJ0&W^VYD\O67
2Z7J\AKT7MLXGN(W+3M?U[5ZPFXX#U]d#J6YBa:<5#EAbP8#H4ENgU+@eD#T/9>A
11(_?TQ18QN,Ua1QdB]H2@REg+U.X=?;5aJ7cTO,R>Q:8B79Gb<AKC>_0VY-1cM2
de:ZG0P#T7H@.;<9(2&[F<A>4E<?GZGFAHW?[)E)7B8&Z5g/G,c,QA](5#>ZPX>_
?NUMBW<cKbYQ7N5_AAF&52LC[4f9</E1^?^CLM_/10-UdUgNMgR3S)C>cd0.a^DG
.B\)&^X-.[D>0T?&/&QL60+TV52cQAR9)=f:0@d43D8OOAPR^QKEU/^,L5;\Y,10
RL(,:T:Fg+1@2,_SB^:dY@Eg_65TgVB;G_>VaAgW(/)DS\KM-)O#AZ:F^FU)BeK&
?Y^#9,O24YE^OL,Kf:0@9-+ODB:fH6/a9=E&F<^(977I]JKfPACd0++3ZZYF_BTc
6FW+?=@)XO2a24^WJ\UCLYCXa5&6(-D<(>X4O^R8b,8-_#01X\]f;)K<fF^OJf-(
0;A<8XM:T>-#QC/Pc\WWdbQ=<^cK&[F2U:1gadW2/+,VAC6RdJ)YNYQ.&FS;Z^cT
+VAA0B5=@,2,E;SU)=8e>9S+T/,1=Fd]T>1;X(dZFb_BVgPOReK0O,I6.e)bU@Wc
[-C+1a#6&AG38KfM\-Y.6][^@QZ]b]K56Ba>I]0.P932^=K#gM36e>O(6K(6QCLC
_dIg3=,[H:3#>4NSKF0dG&&e<^L\a(JP(UQJRXX0OBLP<R\Y<gS=Y;>BZAYOG=-[
FdOTc6#fQW1P@G&3074:>S/B:Sf6.(BfC)P;DFLdEb-J=+&4-BYB[X65SG-^Ib=d
GPB]P72N>[#BY4\X/=X(H2L6M&eYQ[&6cN^S<WD+Y?5HW/5e6OX/7OC_8De0\f@3
7NDedA/(bO8X;93Hg(Y_O),AO3f3M4M2+9+L&A]];U34^9;/bW;[7V.IMZMGNJ[;
INX7a#3?JG^DE&?8UPC<=/9H2TBVJK4aK2[RGYVM6\OPD[F=NP;T5NHRP1bHL-?R
V1FPf&C;E60Ua6E>&5UCC]bFU#6,L@5KJ#;O\:(,+-]&>E[&2P1PVS^XFA;-WX#3
9&T</5N3VJd]BRBL(PD,F@W?N80T:AC.<3DHI=?J</D+#(19W#g(07W>X&egcY?S
(QDUV,2a3\-^B06OWKY&d[ff4IV,_PPN<^EF2Y__3Y_.@>;0537;W<Y7?.GS)R\1
]E27IF2-A&1#&1)aVW<T6KB:[)]O65KS@/.OT3VU(L[RDM3]7bZB0D=cT>_(/?Y@
.Y09D<@\a3^QGKE6L<d^0#]?;>+_DOcJ77#19CEB\ZT+\&O9ge\.)DZBgUK#J3\[
R_/_^J[[Td]2g5N@28J_CRJAOcDNg\[2FMa?)63>+;-4e&:<>;N;LXS4X=Qe8TZS
ZF)dB5G/D?61,&(A>NR)H.2R>#;@Y_21cBAX^5f<<T5.Z+\RG[.)MW6ae/W_8EKQ
IZYb8d(H^)>e@96\]+PZSWGc99YU5g&.@D?R=6P:g&04EE2gF3I>NXLag_N:5Z&d
SP/)5cH9RB>fP<WdUD_T=9._=Xb?GITM:H>TcR:)]L:S/LFZ,6T&/8=[#0DLD2G]
<2NSNHDJ7EcL@^1.44NR93W.^=I<c#M0GJYB.C8^4C00-3_^2R4Q?XUSZ3S2aZff
=Obc:6K\[(.+)UO?6FI[]/FOPe<86RdKT.K>TQ,gA3R3AMfRP7/7KSJ&7OK<?<YZ
fOEPX>ARaDUb__<d)d+?QSBcPNSY:=IM4@Uf[,#RQYFa^3TJDI4?_[@U\5>-XBL;
PLPIHNV^A=_TYH[&]_@-,ZCCKeU\geYXJ_285-EeM(#-M:0G&g<R.b8fDLH?>L1H
014#^TcaaZAf+Kf=T-Y;U;:f5G/<\V47OH-1JJ8>PW+XL-5J&I3QY6IB=,X;E<9b
[b>)ZC==LJX,P0\_(=N3T]<5@7C\P0J?_(7YK/_g\R:6I7\=3B7_TQ0d+5@+R<^R
4cUK-,EK88U###N[1>;eF0c(\),HBUG]C2G39F\U5=?_BdU[fb>ML-OW]=\MQJ>0
-I][EJ+RHOZFFBFX+F3F?T]22@VA))8JU835_Z[3WK_WdMOSEWLPTHUWa[Pd89dS
gA=<PPb,[F8\Tf5_5QT>-BTNA.(HU;:g\66J8+/HJU=-+7,9;8MWX^AB:6,E]EAP
[fHBZ#_C+X@LW>c<cf@6Q2agMf(F#>J6cc09d<)Z>W7GY:HWYMF.2?L7K53PXS_C
GQ0a^c)A]Z#@Q\Z+dXGASBaBddCf5:,<TeTGU3d1I7aKG,K9#23g1Y\OD.3\1OFe
fXBMbOOV^d2^1WL/XaX0#;[/9C@K0d;BK+YLaa(6eYaGP8Z.GaBJAUbVOA&:,C7W
&NJ4A#(6_OVd9/UF[M+Z&V<6H@dMeZF/P&HH([]Y,TYA71Zea1aO9?34^T[B[>M:
,:CD1Ng.3QO30]G5L&HaO3VW+I4Q@=8RE0;.JT:]X@KOa.\K5a1PH0bCeBP\9C4\
;a4X]/3A<]G_@WN^F4DQfc@)Z:M@OP;U#-Aa.W.GaH)(<4Tg5V54;dTHCZT(AYAK
<;Zfb&-10bDWEBF5Q)fP^E1IF]R-Lb[Y^IV?I5D540/e6WP^81c\bT609?OXG&Og
cPfNe&YRIe3[U2Z#6;Odb:<,J^AN/LJ50.8/VGKXDLMdH1OgX42bQ7=JE7<QA;]5
P4[R9]W6>V2IJc3KG;XR0DQ.T8dY\91B7g50/YI&6MJ&Ha@/K>EJ_5UI?QDPH>,S
9N7\<NC\,0B:Y7eAVPK(REZG1-BOc;+DN>J5.2@R=f(<D#PAZ46C27BdDY7?O3&P
LeIbVFG8V,C:+F2_I9-@O=I&T>(E;,J[/aKR@eFP#dHM82XWW,\BPcM.1#2OLP&G
MWF9Aec6,K&2OZW86_+\(9JCE^_g^,gZfV@>028K,FLW/O5J.JKC:cc\KLGV2ROg
Ue4SD<fN67@IFGD5dFDK/.gY#4_OL74SKf>=I,L_PLIIKW8<RD&]fSPZ:Pc])F)D
D1VKK>a.><M#-Hf<)FXO\-RaNOUfL_\:Eg;[;Z(@6#F<9FS;Y1NZ)=&;?LQFPd2H
[E6GH([A[gB^VT5Lda\I<V1)G:)12.,cJZ3[&R8^/fP0eX>DWW5S@a(]c47gWT4Q
&dP@aBeVCc23ZP?G_bCd;DR_,V0PJ<&#TLG^<>aNW7]/<:2-)MGTS&CFdQ@5gQJf
38/8dWZ4ddEZQ3.gMJ<)2V8;MBQ11g0I_I^g.ggW9KSN)X3Cd(V.&]3+QG0##(28
&<>M/4-]Y:9_DU1:13L=WTLB@]TUB4eN:\-OM^FG.\;L:7,.SF_X]A^?P(ZgQ7fD
B&CI(bZ.6A5/R^KTbYLMR#aeI-<HeH2E5fe;G_N&Q-QNQUA@I0KNZ4eGfe6Y)BLa
<P_fc@L=@7K#A&e2N[6,JKP3#_2Z\[V\GLMMC/S<&eWA;4[ab>BU63/-b@?408.a
K.\E?a_HUG9JKJ+-Qd6((EA6X3;a4MEE^a,VQ5P@M-Kc^Sg5_[.FI@ZUP24?>&fQ
RWAX?M#3HUgB:eU/H@Vd+FBTcMA](^KETCZQ/W_Q//-0UgZACdaPB[(.Y(S#V.&=
:UPV#=MaPHQH=K+1?b_KgXPZL-]J.#^P7?J+7S84+cZ4?F<+K+R)C6CEb;1<\(:K
[KZ^3.=0OI_GAEe@48;QBT)QPcHPHQ@\D#Ud=VI2MV[OY3c08.;:QWWPWTQW>465
>([+=f7NeFL;?H6fFG[9UK&K_L+,;:bFCV>37WGdGeO+5NW9dLV5Mb&&Q)?B7c7C
._-_B2):L56GGY1TCO+YM.],U\Ya-XO]\^_2BCKb=1I;EQM+Y(1WHRUfIf)M#?D5
b)^PT^MS]e8_61I8#\E1<d9d-E5,YWIYe>2GG),[N_6,gg/fe@)LJ&Ag4P^JS?J3
g[]2R39UN66;P7K,)WHM+V-)F>]Q(:)+)?B1Gg8I0)dG?-78+_Y6S)7G7A:-GaFB
?5g[SaV1/G+^6T?f2H7E7ERB41DEN\V;B..<DbA9;JFM=L/WeAEW?B.?\1X2&>]1
O8ef(SBVT6Xf_IZ:>fL\Z._<Y=+-3=;B0?afMH,I=RF^=TF]1bOZBMaS#X;L64[>
#(2\5g5+831d8)]9WN0^gegZUQ88[)C5X_8MX0Z)ISVRPD+9?RgT8=4UFb8V8L>1
=(c#YJ@ZRd+121b&5M0OYLV^2[><QR#d4f#WM/LK,[FI@1Q:JdNbX]3d+U04ZSY=
48&gM@/58eH5gIH-OP\BK8@(GCTa2L=NY,.<],K_0#O,Q#>5RQ65O/3g-.6.Q/#e
NRLgQ>1T3.EIcTEE1^8?HLQ32RJSY0C:0[-T.<2gV+WQ>FI2DCCD)(1Z9ZSXc;[S
OA5]b:gbbNCB:)eN-BXFQV>CZCWV2;I2JJ&0U,FRMGAfG5bNfGI^W[?Yf<L/?=94
2Xf-H]=]6c(9+ME^/FLb;3;@Z\.Bc;M4:4<\-YOb<TF9ZP1TG(&c.bO87#C@O#0;
6/<+26.CM2IbYFe,LNcCJ5_Ha72\7(WT>-L:FQg,JZCU5A&IKJ/U,[X2_R,8H]fZ
e/@F=X.Lf)UT=1GTBcQ7M;@4.G)IY8dIb7V:1)0_=_5GWAa,;Y-^BWF_@21XK:VI
<Z-dcKccV>a.__\/-TZ,EKY\cc#gAL-b]56.[e.+K[3[H,032L5XbZ;]B06WFU]W
ZIGJFA0555YR=e0BaWTRMTE@#W@4\6KT8g<&EVaJK:]@Qd]0YD=PT0&Q2@=\3X,,
dZ+B1#5Q9-+P;)Y/AFN8(&F65^U5Y-D\WZ&7ZQ702JIUU.[gBS4J^f1DA;29WLZg
;OJ;84F5,-+3(4dbY5D&1,UL<g)F_1GKge&]SE3>g^FLT=[)42E9P=@Ia0<&0-9f
,D9G1<+FZaE0HO6V+,eWD8G9\dDW>F_=bE[Mg/Z3DE00/LNL:CcXPEFX=.JV5d,-
FL+.>Yd0<>J=5<6\>3Rc;2_X>7(&c]1X@<B@M4>BZJJN,5X?Q+8ge(UR6)Sce7]F
@/&5O+5gQZRHV@+<S5bSKRCd?LKaI]\8@IJI9[YK/Q\9DWJIUN?^E;62-Z+0O>0=
c@XDb4B#Aa3fRNIDPQ_F=0/g);Y(BT;4+KAQgX1EYbL><^27e]G,fGE-,A//9Pg]
T&^^/8N849Mf+dSfg&5NXc6,UC1^e7^/=,9Y4d348C_D,/Z7Z;AL8/TeCIc)c9CE
C/+DSEDO?[H##ccI_I=7:@6BU&Z6MK,0U-3c=ZZO7D9[H2^#WLd5YPMB9LH^PT2g
=AU>#XTWMg7CA?L95Xe)G-eB>f)1M^DW+I&]X0FO;TGG[1Oc>5Ad_]#+(+1dZ^,<
W[\I.LY0<U.?,<,<:ELce]=G2PGOdAA>gK<6J3CN2.S2[4X4,5^R/cdX&?g+cQ&R
-P\4+]=W+(Q/<Y:8/L=L4/]UcD45S(1P/W?H6YU<]e;6(MNXea[&[3TX[/9[U4KE
DPZKe>DA9-E:/V)1cL[1R;W9aD6EMMVRVFPC,EX=+b0AgQ>_\aBI11<PVD6SQa+g
0aPeYO51W@UO;a7+#.CQ?Ae\;ZDE4/M+MDBJ(1]\@QL\^5?#B1J?W)Ya,(MQ1YPg
PC=OGe1E290VG,9>3\).E-g_K1+T)gA,OF8H^QSCFI[DKf6AZf3Y]=EYM6I/L1./
ODc-aD^WB644fc<</2QFJ\^Q9@)7bG]g,1W@K>0<;)[>IJ/L[4gaIG&SZI#dSV28
<&(U[)cKF=/T^0+&K\/PO^-=CG<FEe0.+>#OS@@E<UHT[M].gC@4;7J204O>H\SU
0f2N>F&fCgS)ba3Z=U968-^;UOaAIVL\?J#Xd_48?V<9G&#/[#K^[^BbX/IP0I_X
DB4A=/WQd,dYS/:A;DW;A-PT#U>V@Ld5e=EB]e<\[[=;PYF7B#.IV29O^4(,:Ie#
\I:4E)CEd/N=(>5_(LD,C#I;J=(,NVCaNJTZ8\PYHF..@I\YMBR)?O>,.>ODfIa\
QHD:T9bKGWB??UdT7,GUM2R.[P,_<1[O>d52[YA1S4HZ_VG3,3L9?,&52(GKGL)&
A?^?4M;_9[g(RXO2N6)TfeD59B>BHHMMLVfd>A1G]PE?Q)KbI-9Q4,J:/e_c(#X;
M.g(BNP:(?I/g7?gBYK^M<=P,U9=KXeN6981\AT\ZX9?D)M:KGHQ++UC?U5(UDdb
.H/J89UA?4MN8?cSO\+>#GBQeSd5=5QU>=3)F(7Q_&32PYS1a67_,XBV+K/OR?,H
4O6<b[@N@?[2-KbAIJD\^(g#12YCUODT[1R(cEZ/?4EY.V@Bg2^QFVBS/#=Y/^-D
H5ba\]X#)&K.9]J()gF(<^.;@/5-B>TKb2>Nb8_Z8?Nf4f(/T?6cN8V>>G^G20:-
C)MWQH99J?UAN=W]8D6b@b=07aJU/AMV:+3G@HE?:M25_2(<N9@N)E;>Iag46;G9
LKaB;E]<1U-VWQ&dR\9PYK8)2e26UMF\GGU_/EURE:)FRQKf&Je5@e).N5[G-=XE
O;290g(4a6SLR7D05C<&2&J?O9F625BV+5@7YKTYA5^T3c&C)\ZO>74gb_QM8L_@
M0[#;MN(?181W8RHUD&\00G3M50e4&TANd:^@KAf)X&(=\0Ff2RMDba1UGdZN>&:
?.Edd1L.T\:;a5N_32d\+NSS#T,R7XYB7b8XTAf>WcXP@YP)]E&MXK1UXHY8/7#+
e(Gb<aZ;\.gG1ZP7#Ve;FZIMDZdV7#4<BFd@E)+H8YH22+,IN:HYXR)AI;LY8VeM
6\2[GQ[6Jee6XHL=_]A=Ub4Lf;W_=e/+#ef[CV,+SW#dDADA[<YL(@V+EeBNS0e\
&C3>+)6;?\&g20^>)#dbQ@@>VIEF\e0(A1F&Q=/:Rd&>?RUMIF=[LBRIScCcCGED
9D0ZTA,<\e4H1I\ZK)B\]d+[=bc2a&-LNYX&QW<4(>Z#R9CE;e+;?NJGeML7f>HE
01_eS-_+d([-E)=,_dU1MZ&H8NP&+2(c:@6#dL8#?(Z>aDMCFBP98HAP8:XV&Db8
eJ,9J.OaOIA0Z1g__Z<,cKCH4;ad=dVNWK,EZ^NcUb12d7fROF+^T9A=<M:>#92E
B[(4&ZOd=9BKA008b-R#ZV8\10C:RXQ,gd:?,GLc=GQ@=S.c6g+STP<M66Z+9S+X
c]72QA)P]Lg=9EZ2=ab]5E[CPO0DEK5D\E.b2=H<HVLY/,b)9A]0c=e<&#[Z8I#:
I#Q2BLIXfV,<-\-+4OO,Z\e)QdQ4Bb0Lb6_3[\CNg<WRZEHK^><EL>G3#XA11\2&
&[D@])YIgD_&Z60YY=8:<Q+J(JDY0A[U[F+]U<bU8c>=8X:K3&S@S2KJeO<YZC(@
JZ3DB]5AR<W#\43\>L<aZY+/J0=PfEVb2O75GP+\A69&#;9R]N5GV.KQFb8?85g8
B,6NNK9LTKg>T(D,8EQOICRMJB&13]PMB.EY&eK6g_K>7gVBH651RGDK82MS/<4=
Y=#Y>\eFNF91IB5TEQKI1dNF_dECRb:NZ,AW3^I@Z):Q&(GZ7H^bU6FBI?fRO:4^
^LZXT-\VFLDg\PE)KV=g3J7bfNEa6V?SAEeaNKP<Y[5W>[1>#(S?ba08(WHPGI/8
P\\U7VMIR0,PB:2L>UL\ZDT,S]+dV0\J1WF@ZQJPFOF^;KO34&H[DQfGH4?f@\TF
c#E\I&UPbecJ:8L,b4:&fXQ,)Y@AZ-W=DQGf1>&1O^>QW3IdgG:<QLI\-3;G>#+g
Q-N7J<:,POSUIAa0FZD<?LWdXA?KPa3+\R<Re+;9IAH3:(6af=6D^4\?^D_/5NQE
MP2M9&Qa#79fO]eUT-aGILB(NA,KQEAK4NcFfYC-PZMD^9K+4:B-T0Uc:5.eL<B-
cWAEBCPdB+^?TYZ/;E(6ZfBMfP)AfOABFQ_fSEcT2=:XQSSI4C3bNUKI4We;^UVE
?XgW);H(OO&Xf1^1H:Y3aRGKM>Yf_XNYe6c1<,g8VA[;?]d/fTC]c>ZQ0#TQC\]N
JYT&\\ZAfC92I/62GQ&:,_M\bUM3J=R+bSSG-@2@>>1e)]c(ae1O\R[:fV1c0M<K
bNF5UN910:4@Nf/P>G0<67^Na<I//dc<?&[9?Q7[1_bE3+/K1\E]b1c.G3/f1KB+
^VFG,Y0QeIMQ3d\)\bF]S&g>82>)KGgP0KQPA=OL0FO;YWE05E,NV6U8f(T&VSR)
>caE(c#MTaI7X(30H2W[;<Uf&8^:Ta9e.+bCD(\^Mc:99@/6eWQ7ITAg?6J6d?U7
\KeR9YET1D8OE\bUH1@[13OOLM=H<e(Xb[IFN1KN^YBZI)?6:/[RcBdTIS-^S\^AU$
`endprotected
endmodule